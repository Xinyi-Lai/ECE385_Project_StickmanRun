module digits_rom ( input [7:0] addr, output [7:0] data);

	parameter ROM_LENGTH = 16*10;
	parameter DATA_WIDTH = 8;

	// ROM definition				
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {

		// code x0
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11001110, // 5 **  ***
		8'b11011110, // 6 ** ****
		8'b11110110, // 7 **** **
		8'b11100110, // 8 ***  **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x1
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00011000, // 2
		8'b00111000, // 3
		8'b01111000, // 4    **
		8'b00011000, // 5   ***
		8'b00011000, // 6  ****
		8'b00011000, // 7    **
		8'b00011000, // 8    **
		8'b00011000, // 9    **
		8'b00011000, // a    **
		8'b01111110, // b    **
		8'b00000000, // c    **
		8'b00000000, // d  ******
		8'b00000000, // e
		8'b00000000, // f
		// code x2
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b00000110, // 4      **
		8'b00001100, // 5     **
		8'b00011000, // 6    **
		8'b00110000, // 7   **
		8'b01100000, // 8  **
		8'b11000000, // 9 **
		8'b11000110, // a **   **
		8'b11111110, // b *******
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x3
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b00000110, // 4      **
		8'b00000110, // 5      **
		8'b00111100, // 6   ****
		8'b00000110, // 7      **
		8'b00000110, // 8      **
		8'b00000110, // 9      **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x4
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00001100, // 2     **
		8'b00011100, // 3    ***
		8'b00111100, // 4   ****
		8'b01101100, // 5  ** **
		8'b11001100, // 6 **  **
		8'b11111110, // 7 *******
		8'b00001100, // 8     **
		8'b00001100, // 9     **
		8'b00001100, // a     **
		8'b00011110, // b    ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x5
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111110, // 2 *******
		8'b11000000, // 3 **
		8'b11000000, // 4 **
		8'b11000000, // 5 **
		8'b11111100, // 6 ******
		8'b00000110, // 7      **
		8'b00000110, // 8      **
		8'b00000110, // 9      **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x6
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111000, // 2   ***
		8'b01100000, // 3  **
		8'b11000000, // 4 **
		8'b11000000, // 5 **
		8'b11111100, // 6 ******
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x7
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111110, // 2 *******
		8'b11000110, // 3 **   **
		8'b00000110, // 4      **
		8'b00000110, // 5      **
		8'b00001100, // 6     **
		8'b00011000, // 7    **
		8'b00110000, // 8   **
		8'b00110000, // 9   **
		8'b00110000, // a   **
		8'b00110000, // b   **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x8
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11000110, // 5 **   **
		8'b01111100, // 6  *****
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x9
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11000110, // 5 **   **
		8'b01111110, // 6  ******
		8'b00000110, // 7      **
		8'b00000110, // 8      **
		8'b00000110, // 9      **
		8'b00001100, // a     **
		8'b01111000, // b  ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000 // f
	};

	assign data = ROM[addr];

endmodule  




module stickman_rom ( input [9:0] addr, output [55:0] data);

	//parameter ADDR_WIDTH = 10;
	parameter ROM_LENGTH = 80*9;	// 720
	parameter DATA_WIDTH = 56;
				
	// ROM definition: height: 80*9, width: 56
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {
		// height: 80, width: 56
		//Page 1
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000100000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000011100000000000,
		56'b00000000000000000000000000001111111110000111110000000000,
		56'b00000000000000000000000000011111111000000111110000000000,
		56'b00000000000000000000000011111111100000001111110000000000,
		56'b00000000000000000000011111111111100000001111100000000000,
		56'b00000000000000000001111111111111110000011111100000000000,
		56'b00000000000000001111111111111111111000011111000000000000,
		56'b00000000000000001111111111111111111100111111000000000000,
		56'b00000000000000011111111110011111111100111110000000000000,
		56'b00000000000000011111110000011111111111111110000000000000,
		56'b00000000000000011111000000011111111111111100000000000000,
		56'b00000000000000011111000000011111111111111100000000000000,
		56'b00000000000000011111000000011111011111111000000000000000,
		56'b00000000000000011111000000011111001111111000000000000000,
		56'b00000000000000111110000000011110001111110000000000000000,
		56'b00000000000000111110000000011110000111110000000000000000,
		56'b00000000000000111110000000111110000111100000000000000000,
		56'b00000000000000111110000000111110000001000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111100000000111110000000000000000000000000,
		56'b00000000000001111100000000111110000000000000000000000000,
		56'b00000000000001111100000000111110000000000000000000000000,
		56'b00000000000001111100000000111110000000000000000000000000,
		56'b00000000000000111100000001111110000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111111000000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000011111111111111111110000000000000,
		56'b00000000000000000000000011111111111111111111110000000000,
		56'b00000000000000000000000011111001111111111111111000000000,
		56'b00000000000000000000000111111000000111111111111000000000,
		56'b00000000000000000000000111110000000000011111111000000000,
		56'b00000000000000000000001111110000000000001111110000000000,
		56'b00000000000000000000001111100000000000001111100000000000,
		56'b00000000000000000000001111100000000000011111100000000000,
		56'b00000000000000000000011111100000000000111111000000000000,
		56'b00000000000000000000011111000000000000111111000000000000,
		56'b00000000000000000000111111000000000001111110000000000000,
		56'b00000000000000000000111110000000000001111100000000000000,
		56'b00000000000000000000111110000000000011111100000000000000,
		56'b00000000000000000001111100000000000111111000000000000000,
		56'b00000000000000000011111100000000000111110000000000000000,
		56'b00000000000000000111111100000000001111110000000000000000,
		56'b00000000000000011111111000000000011111100000000000000000,
		56'b00000000000000111111110000000000011111100000000000000000,
		56'b00000000000001111111100000000000011111110000000000000000,
		56'b00000000000011111111000000000000011111110000000000000000,
		56'b00000000000111111100000000000000000111110000000000000000,
		56'b00000000011111111000000000000000000011110000000000000000,
		56'b00000000111111110000000000000000000001100000000000000000,
		56'b00000001111111000000000000000000000000000000000000000000,
		56'b00000011111110000000000000000000000000000000000000000000,
		56'b00000111111100000000000000000000000000000000000000000000,
		56'b00000111111000000000000000000000000000000000000000000000,
		56'b00000011111000000000000000000000000000000000000000000000,
		56'b00000011111000000000000000000000000000000000000000000000,
		56'b00000011111000000000000000000000000000000000000000000000,
		56'b00000001111000000000000000000000000000000000000000000000,
		56'b00000000100000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 2
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000011111000000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100111100000000000,
		56'b00000000000000000000000000111111111111101111100000000000,
		56'b00000000000000000000000000111111111111001111100000000000,
		56'b00000000000000000000000000011111111110001111100000000000,
		56'b00000000000000000000000000001111111100001111100000000000,
		56'b00000000000000000000000000011111110000011111000000000000,
		56'b00000000000000000000000011111111110000011111000000000000,
		56'b00000000000000000000001111111111111000011111000000000000,
		56'b00000000000000000001111111111111111100011111000000000000,
		56'b00000000000000000111111111111111111110111111000000000000,
		56'b00000000000000001111111111111111111111111110000000000000,
		56'b00000000000000001111111110011111111111111110000000000000,
		56'b00000000000000001111111000011111011111111110000000000000,
		56'b00000000000000001111000000011111001111111110000000000000,
		56'b00000000000000011111000000011111000111111110000000000000,
		56'b00000000000000011111000000011111000011111100000000000000,
		56'b00000000000000011111000000011110000001111100000000000000,
		56'b00000000000000011111000000011110000000111000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000111111000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000001111100000000000000000000000000,
		56'b00000000000000011100000001111111100000000000000000000000,
		56'b00000000000000000000000001111111111110000000000000000000,
		56'b00000000000000000000000011111111111111110000000000000000,
		56'b00000000000000000000000011111111111111111111100000000000,
		56'b00000000000000000000000111111111111111111111110000000000,
		56'b00000000000000000000001111110000111111111111111000000000,
		56'b00000000000000000000001111100000000011111111111000000000,
		56'b00000000000000000000011111100000000000001111111000000000,
		56'b00000000000000000000111111000000000000000011111000000000,
		56'b00000000000000000000111110000000000000000111110000000000,
		56'b00000000000000000001111110000000000000000111110000000000,
		56'b00000000000000000011111100000000000000000111110000000000,
		56'b00000000000000000011111100000000000000000111110000000000,
		56'b00000000000000000111111000000000000000000111110000000000,
		56'b00000000000000001111110000000000000000000111110000000000,
		56'b00000000000000011111100000000000000000001111100000000000,
		56'b00000000000001111111100000000000000000001111100000000000,
		56'b00000000000011111111000000000000000000001111100000000000,
		56'b00000000000111111110000000000000000000001111100000000000,
		56'b00000000011111111100000000000000000000001111100000000000,
		56'b00000000111111110000000000000000000000001111100000000000,
		56'b00000011111111100000000000000000000000011111000000000000,
		56'b00000111111110000000000000000000000000011111100000000000,
		56'b00011111111100000000000000000000000000011111110000000000,
		56'b00111111111000000000000000000000000000001111111000000000,
		56'b00111111100000000000000000000000000000000111111000000000,
		56'b00111111000000000000000000000000000000000001110000000000,
		56'b00111110000000000000000000000000000000000000000000000000,
		56'b00111110000000000000000000000000000000000000000000000000,
		56'b00111110000000000000000000000000000000000000000000000000,
		56'b00011110000000000000000000000000000000000000000000000000,
		56'b00001100000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 3
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111000000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111101000000000000000,
		56'b00000000000000000000000001111111111111111100000000000000,
		56'b00000000000000000000000000111111111111111110000000000000,
		56'b00000000000000000000000000111111111111111110000000000000,
		56'b00000000000000000000000000011111111111111110000000000000,
		56'b00000000000000000000000000011111111110111110000000000000,
		56'b00000000000000000000000000001111111100111110000000000000,
		56'b00000000000000000000000000011111110000111110000000000000,
		56'b00000000000000000000000001111111110000111110000000000000,
		56'b00000000000000000000000111111111111000111110000000000000,
		56'b00000000000000000000011111111111111110111110000000000000,
		56'b00000000000000000001111111111111111111111110000000000000,
		56'b00000000000000000011111111111111111111111110000000000000,
		56'b00000000000000001111111111011111011111111110000000000000,
		56'b00000000000000001111111100011111001111111110000000000000,
		56'b00000000000000001111110000011111000111111110000000000000,
		56'b00000000000000001111100000011111000011111110000000000000,
		56'b00000000000000001111100000011111000000111110000000000000,
		56'b00000000000000001111100000011110000000011100000000000000,
		56'b00000000000000000111100000011110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110001111100000000000000000000000000,
		56'b00000000000000000111110001111111100000000000000000000000,
		56'b00000000000000000011100001111111111100000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111111110000000000000,
		56'b00000000000000000000000011111111111111111111100000000000,
		56'b00000000000000000000000011111000011111111111110000000000,
		56'b00000000000000000000000111111000000111111111111000000000,
		56'b00000000000000000000000111110000000000011111111000000000,
		56'b00000000000000000000000111110000000000000011111000000000,
		56'b00000000000000000000001111100000000000000011111000000000,
		56'b00000000000000000000001111100000000000000011111000000000,
		56'b00000000000000000000001111100000000000000011111000000000,
		56'b00000000000000000000011111100000000000000001111000000000,
		56'b00000000000000000000011111000000000000000001111100000000,
		56'b00000000000000000000011111000000000000000001111100000000,
		56'b00000000000000000000111110000000000000000001111100000000,
		56'b00000000000000011111111110000000000000000001111100000000,
		56'b00000000011111111111111110000000000000000001111100000000,
		56'b00001111111111111111111110000000000000000001111100000000,
		56'b00011111111111111111111100000000000000000000111100000000,
		56'b00011111111111111111100000000000000000000000111110000000,
		56'b00111111111111110000000000000000000000000000111110000000,
		56'b00111111000000000000000000000000000000000000111111110000,
		56'b00111110000000000000000000000000000000000000111111110000,
		56'b00111100000000000000000000000000000000000000111111110000,
		56'b00111100000000000000000000000000000000000000011111110000,
		56'b00000000000000000000000000000000000000000000000001000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 4
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000111111111110000000000000000000000,
		56'b00000000000000000000001111111111110000000000000000000000,
		56'b00000000000000000000011111111111110000000000000000000000,
		56'b00000000000000000000111111111111110000000000111000000000,
		56'b00000000000000000000111111011111110000011111111100000000,
		56'b00000000000000000001111110011111111011111111111100000000,
		56'b00000000000000000001111100011111111111111111111100000000,
		56'b00000000000000000001111100111111111111111111111000000000,
		56'b00000000000000000000111100111111111111111111000000000000,
		56'b00000000000000000000111110111111111111110000000000000000,
		56'b00000000000000000000111110111111111100000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111100000000000000000000000000,
		56'b00000000000000000000011111111100000000000000000000000000,
		56'b00000000000000000000011111111110000000000000000000000000,
		56'b00000000000000000000011111111111000000000000000000000000,
		56'b00000000000000000000011111111111100000000000000000000000,
		56'b00000000000000000000011111111111110000000000000000000000,
		56'b00000000000000000000001111111111111000000000000000000000,
		56'b00000000000000000000000001111111111100000000000000000000,
		56'b00000000000000000000000011111011111110000000000000000000,
		56'b00000000000000000000000011111001111111000000000000000000,
		56'b00000000000000000000000011111000111111110000000000000000,
		56'b00000000000000000000000011111000011111111000000000000000,
		56'b00000000000000000000000011111000000111111100000000000000,
		56'b00000000000000000000000011111000000011111110000000000000,
		56'b00000000000000000000000011110000000001111110000000000000,
		56'b00000011111100000000000111110000000000111110000000000000,
		56'b00000111111111111100000111110000000000011111000000000000,
		56'b00001111111111111111111111110000000000011111000000000000,
		56'b00001111111111111111111111110000000000011111100000000000,
		56'b00011111111111111111111111110000000000001111100000000000,
		56'b00001111000001111111111111100000000000001111110000000000,
		56'b00000110000000000011111111100000000000000111110000000000,
		56'b00000000000000000000000111000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000111111000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000001111100000000,
		56'b00000000000000000000000000000000000000000001111100000000,
		56'b00000000000000000000000000000000000000000001111100000000,
		56'b00000000000000000000000000000000000000000000111111110000,
		56'b00000000000000000000000000000000000000000000111111110000,
		56'b00000000000000000000000000000000000000000000111111110000,
		56'b00000000000000000000000000000000000000000000011111110000,
		56'b00000000000000000000000000000000000000000000000010000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 5
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000001111111111000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111111110000000000000000000000,
		56'b00000000000000000000000011111111111111110000000000000000,
		56'b00000000000000000000000011111111111111111111000000000000,
		56'b00000000000000000000000011111111111111111111000000000000,
		56'b00000000000000000000000001111111111111111111000000000000,
		56'b00000000000000000000000001111110011111111111000000000000,
		56'b00000000000000000000000001111110000000000110000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111110000000000000000000000,
		56'b00000000000000000000000001111111111000000000000000000000,
		56'b00000000000000000000000001111111111100000000000000000000,
		56'b00000000000000000000000000111111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111100011111110000000000000000,
		56'b00000000111111000000000000111110011111110000000000000000,
		56'b00000001111111111000000000111110001111111000000000000000,
		56'b00000001111111111110000000111110000111111100000000000000,
		56'b00000001111111111111110000111110000001111110000000000000,
		56'b00000000111111111111111100111110000001111110000000000000,
		56'b00000000000000111111111111111110000000111111000000000000,
		56'b00000000000000001111111111111110000000011111000000000000,
		56'b00000000000000000011111111111110000000011111000000000000,
		56'b00000000000000000000011111111110000000011111100000000000,
		56'b00000000000000000000000011111110000000001111100000000000,
		56'b00000000000000000000000000111100000000001111100000000000,
		56'b00000000000000000000000000000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000011111100000000,
		56'b00000000000000000000000000000000000000000001111111100000,
		56'b00000000000000000000000000000000000000000001111111110000,
		56'b00000000000000000000000000000000000000000001111111110000,
		56'b00000000000000000000000000000000000000000000111111100000,
		56'b00000000000000000000000000000000000000000000011111000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 6
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000011111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000011111111111100000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000001111111111000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000000111111111000000000000000000000,
		56'b00000000000000000000000000111111111100000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111110000000000000000,
		56'b00000000000000000000000001111111111111111000000000000000,
		56'b00000000000000000000000001111101111111111000000000000000,
		56'b00000000000000000000000001111111111111111000000000000000,
		56'b00000000000000000000000001111111111110000000000000000000,
		56'b00000000000000000000000000111111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111110000000000000000000,
		56'b00000000000000000000000000011111111100000000000000000000,
		56'b00000000000000000000000000011111111100000000000000000000,
		56'b00000000000111111110000000011111111110000000000000000000,
		56'b00000000000111111111100000011111111110000000000000000000,
		56'b00000000000111111111111000001111111111000000000000000000,
		56'b00000000000111111111111110001111111111100000000000000000,
		56'b00000000000011111111111111101111111111110000000000000000,
		56'b00000000000000000011111111111111101111110000000000000000,
		56'b00000000000000000000111111111111110111111000000000000000,
		56'b00000000000000000000001111111111110011111000000000000000,
		56'b00000000000000000000000011111111110011111000000000000000,
		56'b00000000000000000000000000111111110011111000000000000000,
		56'b00000000000000000000000000001111110001111100000000000000,
		56'b00000000000000000000000000000001100001111100000000000000,
		56'b00000000000000000000000000000000000001111100000000000000,
		56'b00000000000000000000000000000000000001111110000000000000,
		56'b00000000000000000000000000000000000000111110000000000000,
		56'b00000000000000000000000000000000000000111110000000000000,
		56'b00000000000000000000000000000000000000111111000000000000,
		56'b00000000000000000000000000000000000000011111000000000000,
		56'b00000000000000000000000000000000000000011111000000000000,
		56'b00000000000000000000000000000000000000011111000000000000,
		56'b00000000000000000000000000000000000000001111100000000000,
		56'b00000000000000000000000000000000000000001111111100000000,
		56'b00000000000000000000000000000000000000001111111100000000,
		56'b00000000000000000000000000000000000000000111111100000000,
		56'b00000000000000000000000000000000000000000111111100000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 7
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111000000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000111111111000000000000000000000000,
		56'b00000000000000000000000111111111110000000000000000000000,
		56'b00000000000000000000000111111111111100000000000000000000,
		56'b00000000000000000000000111111111111111100000000000000000,
		56'b00000000000000000000000111111111111111111000000000000000,
		56'b00000000000000000000000111111111111111111111000000000000,
		56'b00000000000000000000000111111110011111111111100000000000,
		56'b00000000000000000000000011111110000011111111100000000000,
		56'b00000000000000000000000011111110000000111111100000000000,
		56'b00000000000000000000000011111100000000000111000000000000,
		56'b00000000000000000000000011111100000000000000000000000000,
		56'b00000000000000000000000011111110000000000000000000000000,
		56'b00000000000000000000000011111110000000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000000111111110000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000001100000011111111100000000000000000000,
		56'b00000000000000000111111111011111111100000000000000000000,
		56'b00000000000000001111111111111111111110000000000000000000,
		56'b00000000000000011111111111111111111111000000000000000000,
		56'b00000000000000011111111111111111111111000000000000000000,
		56'b00000000000000011111001111111111111111100000000000000000,
		56'b00000000000000011110000000111111111111100000000000000000,
		56'b00000000000000000000000000000111111111100000000000000000,
		56'b00000000000000000000000000000111110110000000000000000000,
		56'b00000000000000000000000000000111110000000000000000000000,
		56'b00000000000000000000000000000111110000000000000000000000,
		56'b00000000000000000000000000000111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111000000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000011111110000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000001111110000000000000000000000,

		//Page 8
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111000000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000001111111111111000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000001111111000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000111111111100000000000000000000000,
		56'b00000000000000000000000111111111100000000000000000000000,
		56'b00000000000000000000001111111111100000000000000000000000,
		56'b00000000000000000000011111111111100000000000000000000000,
		56'b00000000000000000000111111011111100000000111110000000000,
		56'b00000000000000000000111111011111100001111111111000000000,
		56'b00000000000000000001111110011111111111111111111000000000,
		56'b00000000000000000001111100011111111111111111110000000000,
		56'b00000000000000000001111100111111111111111111100000000000,
		56'b00000000000000000011111000111111111111111000000000000000,
		56'b00000000000000000011111000111111111110000000000000000000,
		56'b00000000000000000011111000111111100000000000000000000000,
		56'b00000000000000000011111000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110001111110000000000000000000000000,
		56'b00000000000000000111110001111100000000000000000000000000,
		56'b00000000000000001111100001111110000000000000000000000000,
		56'b00000000000000001111100001111111000000000000000000000000,
		56'b00000000000000001111100001111111110000000000000000000000,
		56'b00000000000000001111100001111111111000000000000000000000,
		56'b00000000000000001111000001111111111110000000000000000000,
		56'b00000000000000000000000001111111111111000000000000000000,
		56'b00000000000000000000000001111101111111110000000000000000,
		56'b00000000000000000000000000111100111111111000000000000000,
		56'b00000000000000000000000001111100001111111110000000000000,
		56'b00000000000000000000000000111110000011111111000000000000,
		56'b00000000000000000000000000111111111111111111000000000000,
		56'b00000000000000000000000000111111111111111111000000000000,
		56'b00000000000000000000000011111111111111111111000000000000,
		56'b00000000000000000000000111111111111111111100000000000000,
		56'b00000000000000000000000111111111111110000000000000000000,
		56'b00000000000000000000001111111111000000000000000000000000,
		56'b00000000000000000000001111111110000000000000000000000000,
		56'b00000000000000000000001111111110000000000000000000000000,
		56'b00000000000000000000000111111110000000000000000000000000,
		56'b00000000000000000000000011111110000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000011111000000000000000000000000000,
		56'b00000000000000000000000011111000000000000000000000000000,
		56'b00000000000000000000000111110000000000000000000000000000,
		56'b00000000000000000000000111110000000000000000000000000000,
		56'b00000000000000000000000111110000000000000000000000000000,
		56'b00000000000000000000001111100000000000000000000000000000,
		56'b00000000000000000000001111100000000000000000000000000000,
		56'b00000000000000000000001111100000000000000000000000000000,
		56'b00000000000000000000011111000000000000000000000000000000,
		56'b00000000000000000000011111000000000000000000000000000000,
		56'b00000000000000000000111111100000000000000000000000000000,
		56'b00000000000000000000111111110000000000000000000000000000,
		56'b00000000000000000000111111110000000000000000000000000000,
		56'b00000000000000000000111111110000000000000000000000000000,
		56'b00000000000000000000000111000000000000000000000000000000,

		//Page 9
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000001111111000000000000000000000,
		56'b00000000000000000000000000111111100000000000011000000000,
		56'b00000000000000000000000001111111100000000000111100000000,
		56'b00000000000000000000000111111111110000000001111110000000,
		56'b00000000000000000000011111111111110000000011111100000000,
		56'b00000000000000000001111111111111111000000111111100000000,
		56'b00000000000000000111111111111111111000001111111000000000,
		56'b00000000000000001111111110011111111100011111110000000000,
		56'b00000000000000001111111100011111111100111111100000000000,
		56'b00000000000000001111110000011111111111111111000000000000,
		56'b00000000000000001111100000011111111111111110000000000000,
		56'b00000000000000001111100000011111011111111100000000000000,
		56'b00000000000000001111100000011111011111111000000000000000,
		56'b00000000000000001111100000011110001111110000000000000000,
		56'b00000000000000001111000000111110001111100000000000000000,
		56'b00000000000000001111000000111110000111000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000001111100000000000000000000000000,
		56'b00000000000000011111000001111100000000000000000000000000,
		56'b00000000000000011110000001111111100000000000000000000000,
		56'b00000000000000001100000001111111111100000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111111100000000000000,
		56'b00000000000000000000000001111111111111111111100000000000,
		56'b00000000000000000000000001111100011111111111110000000000,
		56'b00000000000000000000000001111100000011111111110000000000,
		56'b00000000000000000000000001111100000000111111110000000000,
		56'b00000000000000000000000001111000000000111111110000000000,
		56'b00000000000000000000000011111000000001111111000000000000,
		56'b00000000000000000000000011111000000111111110000000000000,
		56'b00000000000000000000000011111000001111111100000000000000,
		56'b00000000000000000000000011111000011111111000000000000000,
		56'b00000000000000000000000011111000111111100000000000000000,
		56'b00000000000000000000000011111011111111000000000000000000,
		56'b00000000000000000000000011111111111110000000000000000000,
		56'b00000000000000000000000011111111111100000000000000000000,
		56'b00000000000000000000000111111111110000000000000000000000,
		56'b00000000000000000000000111111111111000000000000000000000,
		56'b00000000000000000000001111110111111000000000000000000000,
		56'b00000000000000000000011111100011111000000000000000000000,
		56'b00000000000000000000111111000001110000000000000000000000,
		56'b00000000000000000000111111000000000000000000000000000000,
		56'b00000000000000000001111110000000000000000000000000000000,
		56'b00000000000000000011111100000000000000000000000000000000,
		56'b00000000000000000111111000000000000000000000000000000000,
		56'b00000000000000001111111000000000000000000000000000000000,
		56'b00000000000000011111110000000000000000000000000000000000,
		56'b00000000000000011111100000000000000000000000000000000000,
		56'b00000000000000111111000000000000000000000000000000000000,
		56'b00000000000001111110000000000000000000000000000000000000,
		56'b00000000000001111110000000000000000000000000000000000000,
		56'b00000000000001111110000000000000000000000000000000000000,
		56'b00000000000001111111000000000000000000000000000000000000,
		56'b00000000000000111111000000000000000000000000000000000000,
		56'b00000000000000011111000000000000000000000000000000000000,
		56'b00000000000000001110000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000

        };

	assign data = ROM[addr];

endmodule  


module cover_rom ( input [18:0] addr, output [7:0] data);

	//parameter ADDR_WIDTH = 19;
	parameter ROM_LENGTH = 640*480;	// 307200
	parameter DATA_WIDTH = 8;
				
	// ROM definition:
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {
		
		8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 
		8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h83, 8'h7b, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h67, 8'h13, 8'h0, 8'h67, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h42, 8'h0, 8'h0, 8'h5e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h85, 8'h2e, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h67, 8'hd, 8'h0, 8'h1a, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h36, 8'h0, 8'h0, 8'h60, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h87, 8'h29, 8'h0, 8'h0, 8'h6a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h39, 8'h0, 8'h0, 8'h0, 8'h5, 8'he, 8'h27, 8'h5e, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h6b, 8'h2f, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h85, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h81, 8'h64, 8'h48, 8'h3a, 8'h13, 8'h0, 8'h0, 8'h7d, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h8b, 8'h80, 8'h86, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h95, 8'h8d, 8'h6e, 8'h14, 8'h0, 8'h0, 8'h7c, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h7c, 8'h50, 8'h34, 8'he, 8'h1f, 8'h5d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h1a, 8'h0, 8'h0, 8'h13, 8'h83, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h85, 8'h43, 8'h4, 8'h0, 8'h0, 8'h24, 8'hc, 8'h0, 8'h20, 8'h4d, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6e, 8'h0, 8'h0, 8'h5, 8'h69, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h82, 8'h3a, 8'h0, 8'h0, 8'h3, 8'h2e, 8'h65, 8'h48, 8'h16, 8'h0, 8'h0, 8'h2f, 8'h6a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'h35, 8'h25, 8'h54, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h90, 8'h77, 8'h3f, 8'h0, 8'h0, 8'h2c, 8'h62, 8'h89, 8'h94, 8'h8d, 8'h6d, 8'h38, 8'h0, 8'h0, 8'h1a, 8'h5c, 8'h80, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h8b, 8'h8b, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h91, 8'h6f, 8'h2a, 8'h0, 8'h0, 8'h4f, 8'h8e, 8'h95, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h8d, 8'h6a, 8'ha, 8'h0, 8'h0, 8'h36, 8'h81, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h68, 8'h1e, 8'h0, 8'h9, 8'h5e, 8'h8c, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h6d, 8'h23, 8'h0, 8'h0, 8'h12, 8'h6f, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h69, 8'h1e, 8'h0, 8'h14, 8'h63, 8'h8e, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h6e, 8'h32, 8'h0, 8'h0, 8'h6, 8'h47, 8'h82, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h97, 8'h96, 8'h95, 8'h95, 8'h8f, 8'h7c, 8'h72, 8'h84, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h6f, 8'h23, 8'h0, 8'h17, 8'h61, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h79, 8'h46, 8'h8, 8'h0, 8'h0, 8'h2f, 8'h67, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h74, 8'h50, 8'h3a, 8'h37, 8'h37, 8'h37, 8'h37, 8'h33, 8'h1e, 8'h1e, 8'h58, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h88, 8'h65, 8'h29, 8'h0, 8'h15, 8'h5e, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8d, 8'h69, 8'h18, 8'h0, 8'h0, 8'hb, 8'h59, 8'h7f, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h38, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h58, 8'h9, 8'h0, 8'hf, 8'h61, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7f, 8'h39, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h6f, 8'h91, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h62, 8'h9, 8'h0, 8'h38, 8'h37, 8'h3d, 8'h48, 8'h58, 8'h6a, 8'h56, 8'h0, 8'h0, 8'h53, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8e, 8'h4e, 8'h7, 8'h0, 8'h30, 8'h6c, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h4e, 8'h1, 8'h0, 8'h0, 8'h0, 8'h11, 8'h58, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h5a, 8'h6, 8'h10, 8'h84, 8'h84, 8'h86, 8'h89, 8'h8e, 8'h93, 8'h77, 8'h0, 8'h0, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h37, 8'h2, 8'h0, 8'h33, 8'h7a, 8'h92, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h86, 8'h61, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h4f, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5b, 8'h8, 8'h19, 8'h95, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h99, 8'h7b, 8'h0, 8'h0, 8'h3b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h79, 8'h34, 8'h0, 8'h5, 8'h3c, 8'h76, 8'h97, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h82, 8'h4c, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h6c, 8'h96, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h56, 8'h3, 8'h16, 8'h95, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h3b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h74, 8'h2e, 8'h0, 8'h0, 8'h51, 8'h87, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h87, 8'h60, 8'h13, 8'h0, 8'h0, 8'h0, 8'h11, 8'h69, 8'h86, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h4d, 8'h0, 8'h12, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h77, 8'h21, 8'h0, 8'h0, 8'h6a, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h8a, 8'h65, 8'h0, 8'h0, 8'h0, 8'h0, 8'h40, 8'h7f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h4e, 8'h0, 8'h12, 8'h93, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h70, 8'h19, 8'h0, 8'h10, 8'h6d, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h67, 8'h24, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h63, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h59, 8'h4, 8'hd, 8'h8c, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h2c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h61, 8'h18, 8'h0, 8'h1c, 8'h66, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h74, 8'h41, 8'h7, 8'h0, 8'h0, 8'h0, 8'h28, 8'h4f, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h5d, 8'h3, 8'h6, 8'h7a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h0, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h5d, 8'h15, 8'h0, 8'h21, 8'h65, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h89, 8'h62, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h74, 8'h93, 8'h9b, 8'h95, 8'h67, 8'h6, 8'h0, 8'h51, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7c, 8'h0, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h5f, 8'h18, 8'h0, 8'h25, 8'h70, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h79, 8'h37, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h6a, 8'h8a, 8'h97, 8'h78, 8'hb, 8'h0, 8'h18, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7d, 8'h2, 8'h0, 8'h20, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5e, 8'hb, 8'h0, 8'h1f, 8'h7e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h90, 8'h7f, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h93, 8'h81, 8'hf, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7f, 8'hd, 8'h0, 8'h12, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h85, 8'h46, 8'h4, 8'h0, 8'h26, 8'h78, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h5c, 8'h25, 8'h0, 8'h0, 8'h0, 8'h36, 8'h65, 8'hc, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h88, 8'h31, 8'h0, 8'hb, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7d, 8'h42, 8'h0, 8'h5, 8'h34, 8'h6f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h91, 8'h72, 8'h32, 8'h0, 8'h0, 8'h0, 8'h6, 8'h0, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h49, 8'h0, 8'h8, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h77, 8'h3b, 8'h0, 8'h2, 8'h40, 8'h79, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h7a, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h52, 8'h0, 8'h7, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h79, 8'h34, 8'h0, 8'h0, 8'h4c, 8'h82, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h8a, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h81, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h53, 8'h0, 8'h7, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h23, 8'h0, 8'h0, 8'h56, 8'h8b, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h68, 8'h0, 8'h0, 8'h0, 8'h0, 8'h75, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h54, 8'h0, 8'h7, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7c, 8'h2d, 8'h0, 8'hb, 8'h55, 8'h8a, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h53, 8'h0, 8'h0, 8'h0, 8'hd, 8'h6f, 8'h9a, 8'h9b, 8'h9a, 8'h90, 8'h55, 8'h2, 8'h2, 8'h89, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h73, 8'h2d, 8'h0, 8'h4, 8'h4a, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h38, 8'h0, 8'h0, 8'h0, 8'h46, 8'h8b, 8'h9b, 8'h9b, 8'h90, 8'h51, 8'h0, 8'h0, 8'h7c, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h6e, 8'h29, 8'h0, 8'h0, 8'h42, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h75, 8'h2c, 8'h0, 8'h0, 8'h3b, 8'h83, 8'h9b, 8'h9b, 8'h8d, 8'h4b, 8'h0, 8'h0, 8'h73, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h72, 8'h1b, 8'h0, 8'h0, 8'h4c, 8'h83, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h74, 8'h32, 8'h3, 8'h59, 8'h8f, 8'h9b, 8'h9b, 8'h8d, 8'h49, 8'h0, 8'h0, 8'h5f, 8'h84, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h75, 8'h9, 8'h0, 8'h4, 8'h5f, 8'h8b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h96, 8'h87, 8'h7e, 8'h8f, 8'h99, 8'h9b, 8'h9a, 8'h8f, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h76, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h65, 8'h7, 8'h0, 8'h18, 8'h62, 8'h8d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h5f, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8b, 8'h5b, 8'hf, 8'h0, 8'h1b, 8'h64, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h79, 8'h33, 8'h9, 8'h2c, 8'hc, 8'h0, 8'h8, 8'h4d, 8'h81, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h5b, 8'h12, 8'h0, 8'h14, 8'h6d, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h73, 8'h68, 8'h89, 8'h65, 8'h1c, 8'h0, 8'h0, 8'h3e, 8'h76, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h5e, 8'h8, 8'h0, 8'h1d, 8'h80, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h96, 8'h9a, 8'h95, 8'h7e, 8'h3b, 8'h0, 8'h0, 8'h33, 8'h73, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h57, 8'h0, 8'h0, 8'h31, 8'h80, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h47, 8'h0, 8'h0, 8'h12, 8'h5d, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h7f, 8'h46, 8'h0, 8'h0, 8'h39, 8'h78, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h49, 8'h0, 8'h0, 8'h0, 8'h30, 8'h77, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h7c, 8'h43, 8'h5, 8'h0, 8'h3e, 8'h7a, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h4e, 8'h23, 8'h0, 8'h0, 8'h24, 8'h5e, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h87, 8'h4b, 8'hb, 8'h0, 8'h44, 8'h82, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h83, 8'h4c, 8'h0, 8'h0, 8'h10, 8'h53, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h65, 8'hd, 8'ha, 8'h54, 8'h90, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h64, 8'hf, 8'h0, 8'h0, 8'h4e, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h77, 8'ha, 8'h0, 8'h40, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h6e, 8'h25, 8'h0, 8'h16, 8'h79, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h6f, 8'h1b, 8'h0, 8'h38, 8'h7b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h92, 8'h66, 8'h14, 8'hf, 8'h67, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h78, 8'h34, 8'h0, 8'h2b, 8'h73, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h6e, 8'h54, 8'h52, 8'h44, 8'h10, 8'h8, 8'h4b, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8c, 8'h4e, 8'hb, 8'h14, 8'h78, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h79, 8'h68, 8'h48, 8'h16, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h84, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h7c, 8'h2d, 8'h15, 8'h7e, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h69, 8'h9, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h73, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h4f, 8'h23, 8'h3f, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h76, 8'h6c, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7c, 8'h32, 8'h0, 8'h0, 8'h0, 8'hc, 8'h48, 8'h55, 8'h56, 8'h57, 8'h59, 8'h6a, 8'h8e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h67, 8'h56, 8'h6d, 8'h94, 8'h8f, 8'h90, 8'h89, 8'h71, 8'h47, 8'h28, 8'h18, 8'h8, 8'hc, 8'h46, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h89, 8'h71, 8'h59, 8'h4b, 8'h45, 8'h3b, 8'h31, 8'h2c, 8'h33, 8'h47, 8'h61, 8'h74, 8'h76, 8'h74, 8'h71, 8'h6c, 8'h5c, 8'h3c, 8'h3b, 8'h70, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h39, 8'h0, 8'h18, 8'h42, 8'h66, 8'h8a, 8'h94, 8'h92, 8'h93, 8'h94, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h78, 8'h53, 8'h46, 8'h56, 8'h74, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7d, 8'h57, 8'h41, 8'h43, 8'h3e, 8'h3c, 8'h35, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h7c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7b, 8'h46, 8'h13, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h1a, 8'h1d, 8'h1a, 8'h17, 8'h12, 8'h0, 8'h0, 8'h0, 8'h16, 8'h46, 8'h60, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h4a, 8'h0, 8'h62, 8'h8e, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h34, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h65, 8'h82, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6e, 8'h28, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h19, 8'h6, 8'h2c, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'ha, 8'h83, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4d, 8'h0, 8'h6a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h75, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h6b, 8'h96, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h56, 8'h29, 8'h35, 8'h74, 8'h7e, 8'h80, 8'h7e, 8'h80, 8'h6e, 8'h15, 8'h0, 8'h28, 8'h7f, 8'h87, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h37, 8'h0, 8'h0, 8'h1e, 8'h22, 8'h1d, 8'h18, 8'h12, 8'he, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h86, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h4f, 8'h0, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6e, 8'h0, 8'hd, 8'h3b, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h20, 8'h58, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h85, 8'h78, 8'h7f, 8'h95, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h81, 8'h16, 8'h0, 8'h2d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h3f, 8'h0, 8'h0, 8'h5b, 8'h74, 8'h79, 8'h76, 8'h74, 8'h73, 8'h70, 8'h6a, 8'h63, 8'h5f, 8'h60, 8'h5f, 8'h61, 8'h62, 8'h58, 8'h28, 8'h0, 8'h0, 8'h2b, 8'h71, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h4e, 8'h0, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h6b, 8'h0, 8'h34, 8'h7a, 8'h7b, 8'h49, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h34, 8'h5f, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h16, 8'h0, 8'h2e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h3d, 8'h0, 8'h0, 8'h68, 8'h91, 8'h98, 8'h98, 8'h98, 8'h98, 8'h97, 8'h97, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h95, 8'h8a, 8'h53, 8'h0, 8'h0, 8'h4a, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4d, 8'h0, 8'h73, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h66, 8'h0, 8'h35, 8'h85, 8'h98, 8'h92, 8'h7d, 8'h45, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2, 8'h42, 8'h5d, 8'h7c, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h1b, 8'h0, 8'h2f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h39, 8'h0, 8'h0, 8'h63, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h63, 8'h0, 8'h0, 8'h3b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4d, 8'h0, 8'h73, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h5c, 8'h0, 8'h2f, 8'h80, 8'h9b, 8'h9a, 8'h9a, 8'h91, 8'h8a, 8'h7e, 8'h5a, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h65, 8'h7e, 8'h88, 8'h80, 8'h88, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h21, 8'h0, 8'h2a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h3c, 8'h0, 8'h0, 8'h5d, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h71, 8'h0, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4d, 8'h0, 8'h72, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h86, 8'h7e, 8'h7b, 8'h7f, 8'h8d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h91, 8'h55, 8'h0, 8'h26, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h87, 8'h76, 8'h43, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'hd, 8'h2c, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h35, 8'h0, 8'h1f, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h45, 8'h0, 8'h0, 8'h57, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h75, 8'h0, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4d, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h62, 8'h26, 8'h0, 8'h0, 8'h4, 8'h4b, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h53, 8'h0, 8'h24, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h65, 8'h47, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h5c, 8'h0, 8'h13, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h50, 8'h0, 8'h0, 8'h3f, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'h0, 8'h0, 8'h1f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h4a, 8'h0, 8'h70, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h32, 8'h7a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h62, 8'h30, 8'h10, 8'h8, 8'h11, 8'h39, 8'h70, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h86, 8'h40, 8'h0, 8'h20, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h8e, 8'h72, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h71, 8'h6, 8'h7, 8'h6d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h66, 8'h2, 8'h0, 8'h18, 8'h87, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7d, 8'h3, 8'h0, 8'h15, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h49, 8'h0, 8'h6f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h5d, 8'h0, 8'hc, 8'h2e, 8'h42, 8'h4d, 8'h3b, 8'h27, 8'h6, 8'h0, 8'h1b, 8'h4a, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h80, 8'h52, 8'h2f, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h29, 8'h44, 8'h77, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h72, 8'h1c, 8'h0, 8'h17, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8d, 8'h53, 8'h0, 8'h0, 8'h0, 8'hf, 8'h67, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h74, 8'h5, 8'h0, 8'h54, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h79, 8'hc, 8'h0, 8'h0, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h1f, 8'h0, 8'h7, 8'h73, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h48, 8'h0, 8'h6e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h74, 8'h25, 8'h0, 8'h4d, 8'h87, 8'h92, 8'h92, 8'h8e, 8'h82, 8'h53, 8'h16, 8'h0, 8'h0, 8'h41, 8'h81, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h8c, 8'h69, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h69, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h5b, 8'h0, 8'h0, 8'h11, 8'h6b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h85, 8'h24, 8'h0, 8'h0, 8'h2, 8'h66, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h77, 8'h1, 8'h0, 8'h31, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h12, 8'h0, 8'h0, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h37, 8'h0, 8'h0, 8'h5f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9a, 8'h98, 8'h93, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h47, 8'h0, 8'h6d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h4f, 8'h0, 8'h1d, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h80, 8'h4f, 8'h0, 8'h0, 8'h44, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8b, 8'h5d, 8'h9, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h5d, 8'h81, 8'h86, 8'h7f, 8'h5d, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h9, 8'h5c, 8'h8f, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h4a, 8'h0, 8'h0, 8'h18, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h65, 8'h24, 8'h3, 8'h3d, 8'h7d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h1, 8'h0, 8'h12, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h13, 8'h0, 8'h0, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h4b, 8'h0, 8'h0, 8'h46, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h98, 8'h95, 8'h95, 8'h93, 8'h93, 8'h93, 8'h88, 8'h66, 8'h66, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8d, 8'h44, 8'h0, 8'h6a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h45, 8'h0, 8'h58, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h4c, 8'h0, 8'h3, 8'h5c, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h8a, 8'h4c, 8'h0, 8'h0, 8'h0, 8'he, 8'h65, 8'h78, 8'h84, 8'h92, 8'h9a, 8'h9b, 8'h99, 8'h93, 8'h83, 8'h70, 8'h46, 8'h0, 8'h0, 8'h0, 8'h55, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h44, 8'h0, 8'h0, 8'h27, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h32, 8'h0, 8'h0, 8'h0, 8'h9, 8'h13, 8'h20, 8'h36, 8'h6c, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6f, 8'h39, 8'h26, 8'h3e, 8'h75, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h5, 8'h0, 8'h9, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h13, 8'h0, 8'h0, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h63, 8'h0, 8'h0, 8'h1f, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7f, 8'h39, 8'h40, 8'h39, 8'h11, 8'h5, 8'h2, 8'h0, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h41, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h44, 8'h0, 8'h6a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h7f, 8'h57, 8'h2a, 8'h12, 8'h9, 8'h7, 8'h6, 8'h11, 8'h32, 8'h61, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h84, 8'h36, 8'h0, 8'h71, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'h34, 8'h0, 8'h1b, 8'h8b, 8'h9a, 8'h91, 8'h62, 8'h14, 8'h0, 8'h0, 8'h7, 8'h48, 8'h6e, 8'h93, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h85, 8'h57, 8'hc, 8'h0, 8'h0, 8'h6a, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h80, 8'h31, 8'h0, 8'h0, 8'h3a, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h61, 8'h22, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h30, 8'h58, 8'h85, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h83, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h43, 8'h60, 8'h82, 8'h96, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h80, 8'hd, 8'h0, 8'h6, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h46, 8'h0, 8'h0, 8'h0, 8'h29, 8'h46, 8'h4d, 8'h4e, 8'h49, 8'h43, 8'h3f, 8'h44, 8'h53, 8'h6b, 8'h74, 8'h75, 8'h6f, 8'h69, 8'h64, 8'h45, 8'h0, 8'h0, 8'h2, 8'h8d, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8d, 8'h57, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h43, 8'h0, 8'h6a, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h5e, 8'h3b, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h35, 8'h4c, 8'h7f, 8'h97, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h74, 8'h29, 8'h0, 8'h7c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h68, 8'h18, 8'h0, 8'h49, 8'h79, 8'h55, 8'h9, 8'h0, 8'h0, 8'h22, 8'h5e, 8'h8c, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h5a, 8'h5, 8'h0, 8'h24, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h63, 8'h11, 8'h0, 8'h0, 8'h4b, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h88, 8'h74, 8'h4c, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h5a, 8'h6e, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h69, 8'h18, 8'h0, 8'h1a, 8'h8, 8'h0, 8'h0, 8'hd, 8'h3c, 8'h54, 8'h5f, 8'h62, 8'h69, 8'h72, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h13, 8'h0, 8'h4, 8'h92, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h83, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h22, 8'h22, 8'h1a, 8'h11, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h81, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'hd, 8'h10, 8'h11, 8'h14, 8'h13, 8'h0, 8'h0, 8'h4, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h43, 8'h0, 8'h6a, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h7d, 8'h48, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h56, 8'h69, 8'h83, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5f, 8'h17, 8'h5, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8a, 8'h42, 8'h0, 8'h0, 8'h31, 8'h3, 8'h0, 8'h0, 8'h45, 8'h7c, 8'h96, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h8d, 8'h54, 8'h0, 8'h0, 8'h43, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h55, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h92, 8'h8c, 8'h88, 8'h83, 8'h72, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h52, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h4b, 8'h6, 8'hd, 8'h82, 8'h7f, 8'h4e, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h59, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h17, 8'h0, 8'h1, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h62, 8'h90, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'h2c, 8'h0, 8'h0, 8'h27, 8'h7e, 8'h86, 8'h89, 8'h8a, 8'h89, 8'h8a, 8'h8b, 8'h72, 8'h9, 8'h0, 8'h0, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h43, 8'h0, 8'h6a, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h78, 8'h33, 8'h0, 8'h0, 8'h0, 8'h28, 8'h70, 8'h7e, 8'h85, 8'h86, 8'h86, 8'h86, 8'h82, 8'h65, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h79, 8'h90, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h45, 8'h1, 8'h23, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h67, 8'h13, 8'h0, 8'h0, 8'h0, 8'h7, 8'h61, 8'h8c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h48, 8'h0, 8'h11, 8'h64, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8a, 8'h77, 8'h5f, 8'h39, 8'h6, 8'h0, 8'h27, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h34, 8'h0, 8'h1f, 8'h91, 8'h99, 8'h8d, 8'h7f, 8'h71, 8'h65, 8'h51, 8'h3a, 8'h1d, 8'h1, 8'h0, 8'h13, 8'h5c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h1b, 8'h0, 8'h1, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h89, 8'h6d, 8'h46, 8'h2d, 8'h4e, 8'h47, 8'h43, 8'h45, 8'h4b, 8'h4d, 8'h4d, 8'h40, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h10, 8'h5, 8'h0, 8'h0, 8'h0, 8'h78, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h38, 8'h0, 8'h0, 8'h53, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hf, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h44, 8'h0, 8'h6a, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h74, 8'h26, 8'h0, 8'h0, 8'h46, 8'h6f, 8'h83, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h92, 8'h83, 8'h72, 8'h60, 8'h29, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h7d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3c, 8'he, 8'h57, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7d, 8'h32, 8'h0, 8'h0, 8'h19, 8'h6c, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h79, 8'hf, 8'h0, 8'h34, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h24, 8'h0, 8'h0, 8'h0, 8'h60, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h91, 8'h80, 8'h64, 8'h4d, 8'h40, 8'h47, 8'h62, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h25, 8'h0, 8'h3b, 8'h93, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h93, 8'h89, 8'h7d, 8'h6c, 8'h42, 8'h0, 8'h0, 8'h52, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h2f, 8'h0, 8'h0, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h87, 8'h7b, 8'h8a, 8'h87, 8'h84, 8'h87, 8'h88, 8'h89, 8'h89, 8'h83, 8'h75, 8'h64, 8'h5d, 8'h5f, 8'h64, 8'h67, 8'h6c, 8'h68, 8'h4e, 8'h37, 8'h47, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h83, 8'h3a, 8'h0, 8'h1, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'hf, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h41, 8'h0, 8'h67, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h86, 8'h30, 8'h0, 8'h0, 8'h54, 8'h85, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h99, 8'h91, 8'h78, 8'h58, 8'h3d, 8'h14, 8'h0, 8'h0, 8'h0, 8'h31, 8'h79, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h89, 8'h6a, 8'h4b, 8'h34, 8'h2f, 8'h38, 8'h40, 8'h4a, 8'h58, 8'h6f, 8'h8c, 8'h86, 8'h3a, 8'h14, 8'h68, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h88, 8'h41, 8'h0, 8'h0, 8'h55, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h52, 8'h0, 8'he, 8'h74, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h1f, 8'h0, 8'h0, 8'h5, 8'h6c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h89, 8'h56, 8'h35, 8'h17, 8'h1c, 8'h5b, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h1d, 8'ha, 8'h63, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h5c, 8'h16, 8'h0, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h4c, 8'h0, 8'h0, 8'h86, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h9a, 8'h99, 8'h9a, 8'h99, 8'h9a, 8'h99, 8'h99, 8'h99, 8'h96, 8'h96, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h95, 8'h90, 8'h88, 8'h86, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h39, 8'h0, 8'h0, 8'h59, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hf, 8'h0, 8'h0, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h3d, 8'h0, 8'h64, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h42, 8'h0, 8'h5, 8'h54, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h93, 8'h8b, 8'h6c, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h61, 8'h3e, 8'h33, 8'h26, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h16, 8'h31, 8'h40, 8'h1d, 8'h1b, 8'h78, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h57, 8'h0, 8'h40, 8'h80, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h7b, 8'h11, 8'h0, 8'h4c, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h81, 8'h1a, 8'h0, 8'h0, 8'h20, 8'h76, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h78, 8'h5f, 8'h45, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h7e, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h79, 8'h18, 8'h1e, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h65, 8'he, 8'h0, 8'h0, 8'hc, 8'h63, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6a, 8'h10, 8'h0, 8'h77, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h3f, 8'h0, 8'h0, 8'h4f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'hf, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h3b, 8'h0, 8'h62, 8'h93, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h91, 8'h8b, 8'h84, 8'h7b, 8'h73, 8'h70, 8'h74, 8'h7f, 8'h8d, 8'h97, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h68, 8'h0, 8'h0, 8'h48, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h92, 8'h95, 8'h97, 8'h97, 8'h96, 8'h87, 8'h51, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h77, 8'h4d, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h89, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h83, 8'h4e, 8'he, 8'h4a, 8'h6e, 8'h80, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h1d, 8'h0, 8'h2f, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h11, 8'h0, 8'h0, 8'h38, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h73, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h8c, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h65, 8'h10, 8'h2a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8b, 8'h36, 8'h0, 8'h0, 8'h0, 8'h30, 8'h7c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h77, 8'h1d, 8'h0, 8'h6b, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h53, 8'h0, 8'h0, 8'h3b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'hf, 8'h0, 8'h0, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h3a, 8'h0, 8'h61, 8'h92, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h6b, 8'h55, 8'h3e, 8'h1f, 8'h2, 8'h0, 8'ha, 8'h2d, 8'h5a, 8'h80, 8'h8b, 8'h92, 8'h95, 8'h7d, 8'h34, 8'h0, 8'h45, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h84, 8'h6d, 8'h7a, 8'h7e, 8'h8a, 8'h96, 8'h99, 8'h85, 8'h33, 8'h0, 8'h0, 8'h10, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h69, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h66, 8'h7f, 8'h86, 8'h86, 8'h87, 8'h87, 8'h87, 8'h86, 8'h7e, 8'h51, 8'h0, 8'h0, 8'h7, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h84, 8'h4e, 8'h6, 8'h0, 8'h0, 8'h0, 8'h30, 8'h6a, 8'h8b, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h25, 8'h0, 8'h1f, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h86, 8'h85, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5e, 8'h3, 8'h0, 8'h0, 8'h52, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h59, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h48, 8'h6, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7c, 8'h4b, 8'h1, 8'h0, 8'h0, 8'h2f, 8'h7d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7e, 8'h22, 8'h0, 8'h5c, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h68, 8'h0, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h10, 8'h0, 8'h0, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h3a, 8'h0, 8'h62, 8'h93, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h62, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h75, 8'h5c, 8'h0, 8'h10, 8'h66, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7c, 8'h34, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h5c, 8'h9b, 8'h97, 8'h73, 8'h10, 8'h0, 8'h0, 8'h71, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h48, 8'h0, 8'h0, 8'h0, 8'h30, 8'h64, 8'h6e, 8'h82, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8c, 8'h64, 8'hc, 8'h0, 8'h2e, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h6e, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h86, 8'h29, 8'h0, 8'h19, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h65, 8'h18, 8'h0, 8'h34, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h68, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h76, 8'h4a, 8'ha, 8'h0, 8'h0, 8'h27, 8'h69, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h1a, 8'h0, 8'h18, 8'h51, 8'h6b, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h87, 8'h5f, 8'h1b, 8'h0, 8'h0, 8'h10, 8'h48, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h83, 8'h25, 8'h0, 8'h3f, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h71, 8'h0, 8'h0, 8'h23, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h1b, 8'h0, 8'h0, 8'h75, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h3b, 8'h0, 8'h62, 8'h93, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5f, 8'h2c, 8'h21, 8'h34, 8'h3a, 8'h3c, 8'h3c, 8'h3c, 8'h3c, 8'h3a, 8'h32, 8'h1e, 8'h0, 8'h0, 8'h0, 8'h1, 8'h4, 8'h0, 8'h44, 8'h81, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h5a, 8'h1, 8'h0, 8'h4, 8'h1f, 8'hd, 8'h12, 8'h60, 8'h91, 8'h8a, 8'h39, 8'h0, 8'h0, 8'h33, 8'h7c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h8e, 8'h48, 8'h0, 8'h0, 8'h12, 8'h4a, 8'h7d, 8'h94, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h87, 8'h39, 8'h0, 8'hb, 8'h7a, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h50, 8'h0, 8'h0, 8'h41, 8'h52, 8'h51, 8'h4b, 8'h3e, 8'h25, 8'h0, 8'h14, 8'h46, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h21, 8'h0, 8'h26, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h6d, 8'h2e, 8'h27, 8'ha, 8'h0, 8'h33, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h57, 8'h86, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h8c, 8'h5a, 8'h0, 8'h0, 8'h0, 8'hd, 8'h38, 8'h50, 8'h80, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h87, 8'h6b, 8'h64, 8'h74, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h68, 8'h0, 8'h0, 8'h0, 8'h9, 8'h57, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h6c, 8'h19, 8'h0, 8'h0, 8'h0, 8'h34, 8'h65, 8'h89, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h29, 8'h0, 8'h16, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h75, 8'h0, 8'h0, 8'h1c, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h2b, 8'h0, 8'h0, 8'h64, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h3e, 8'h0, 8'h59, 8'h8f, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h7d, 8'h24, 8'h0, 8'h0, 8'h77, 8'h8c, 8'h90, 8'h91, 8'h90, 8'h91, 8'h91, 8'h88, 8'h75, 8'h4b, 8'h13, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h72, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8a, 8'h37, 8'h0, 8'h0, 8'h39, 8'h61, 8'h27, 8'h0, 8'h25, 8'h88, 8'h94, 8'h65, 8'h9, 8'h0, 8'h0, 8'h61, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h71, 8'h10, 8'h0, 8'hb, 8'h65, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h67, 8'h37, 8'h3d, 8'h83, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7f, 8'h1c, 8'h4, 8'h3e, 8'h8f, 8'h93, 8'h94, 8'h92, 8'h8e, 8'h76, 8'h3a, 8'h1d, 8'h16, 8'h46, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h80, 8'h1a, 8'h0, 8'h49, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h73, 8'h30, 8'h36, 8'h61, 8'h53, 8'h8, 8'h0, 8'h31, 8'h65, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h38, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h5c, 8'h75, 8'h80, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8b, 8'h5a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h38, 8'h61, 8'h7e, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h81, 8'h4a, 8'h17, 8'hc, 8'h26, 8'h52, 8'h68, 8'h72, 8'h80, 8'h8f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8e, 8'h56, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6e, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h6d, 8'h21, 8'h0, 8'h0, 8'h0, 8'ha, 8'h49, 8'h78, 8'h93, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h2d, 8'h0, 8'h0, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h79, 8'h0, 8'h0, 8'he, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h45, 8'h0, 8'h0, 8'h41, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h44, 8'h0, 8'h48, 8'h86, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h52, 8'h0, 8'h0, 8'h1b, 8'h8a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h92, 8'h7c, 8'h3a, 8'h5, 8'he, 8'h59, 8'h8b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'h19, 8'h0, 8'h0, 8'h64, 8'h82, 8'h4f, 8'h2, 8'h5, 8'h81, 8'h9a, 8'h89, 8'h3a, 8'h0, 8'h0, 8'h4b, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h43, 8'h0, 8'h0, 8'h55, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h92, 8'h8b, 8'h8e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h59, 8'h0, 8'h27, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8b, 8'h6a, 8'h1d, 8'h19, 8'h7f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h75, 8'h12, 8'h13, 8'h77, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7f, 8'h41, 8'hc, 8'h69, 8'h90, 8'h8e, 8'h5c, 8'h0, 8'h0, 8'h9, 8'h4a, 8'h7f, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h25, 8'h2f, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h94, 8'h7f, 8'h54, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h6c, 8'h90, 8'h96, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h57, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h5e, 8'h82, 8'h91, 8'h92, 8'h93, 8'h95, 8'h94, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h61, 8'h0, 8'h0, 8'h0, 8'h32, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h88, 8'h63, 8'h1a, 8'h0, 8'h0, 8'h0, 8'ha, 8'h74, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h30, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h19, 8'h0, 8'h0, 8'h67, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h68, 8'hf, 8'h0, 8'h4, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h49, 8'h0, 8'h3b, 8'h7e, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7b, 8'h1, 8'h0, 8'h6, 8'h79, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h89, 8'h87, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h74, 8'h8, 8'h0, 8'h0, 8'h7c, 8'h94, 8'h76, 8'h28, 8'h0, 8'h7c, 8'h9b, 8'h92, 8'h54, 8'h0, 8'h0, 8'h35, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h77, 8'h0, 8'h0, 8'h33, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h69, 8'h8, 8'h1, 8'h55, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h84, 8'h2b, 8'h7, 8'h5b, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h56, 8'ha, 8'h2b, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h44, 8'h5, 8'h30, 8'h83, 8'h99, 8'h9a, 8'h89, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h27, 8'h8b, 8'h99, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h41, 8'h5a, 8'h22, 8'h1d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h8c, 8'h75, 8'h58, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h7a, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4c, 8'h0, 8'h1f, 8'h4e, 8'h56, 8'h3d, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h18, 8'h34, 8'h6b, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h44, 8'h0, 8'h13, 8'h7d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h78, 8'h4d, 8'h2, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h7c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h32, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h2b, 8'h0, 8'h0, 8'h57, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h80, 8'h27, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h49, 8'h0, 8'h35, 8'h7d, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h61, 8'h0, 8'h0, 8'h22, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h5e, 8'h0, 8'h0, 8'h1, 8'h85, 8'h9a, 8'h8a, 8'h3c, 8'h0, 8'h6a, 8'h93, 8'h96, 8'h73, 8'h1b, 8'h0, 8'h5, 8'h60, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h4c, 8'h0, 8'h26, 8'h78, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6a, 8'h1f, 8'h59, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h2a, 8'h7, 8'h60, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h1d, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h46, 8'ha, 8'h1a, 8'h7b, 8'h95, 8'h9b, 8'h9b, 8'h98, 8'h8a, 8'h5c, 8'h1b, 8'h0, 8'h0, 8'h25, 8'h71, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h4e, 8'h0, 8'h0, 8'h2f, 8'h72, 8'h49, 8'hb, 8'h1e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h79, 8'h43, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9, 8'h31, 8'h5f, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h90, 8'h48, 8'h0, 8'h45, 8'h82, 8'h90, 8'h84, 8'h67, 8'h45, 8'h30, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h5d, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h86, 8'h2e, 8'h0, 8'h29, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8a, 8'h60, 8'h32, 8'h0, 8'h0, 8'h0, 8'h32, 8'h70, 8'h77, 8'h51, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h45, 8'h0, 8'h0, 8'h6b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h35, 8'h0, 8'h0, 8'h53, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h33, 8'h0, 8'h0, 8'h5d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h47, 8'h0, 8'h2c, 8'h7a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h27, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8b, 8'h41, 8'h0, 8'h0, 8'h20, 8'h89, 8'h9b, 8'h8f, 8'h40, 8'h0, 8'h54, 8'h8a, 8'h98, 8'h87, 8'h46, 8'h0, 8'h0, 8'h4a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h74, 8'h20, 8'h0, 8'h48, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h68, 8'h8a, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h25, 8'ha, 8'h6f, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h6c, 8'h2, 8'h1f, 8'h6b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h46, 8'he, 8'h1e, 8'h65, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h6f, 8'h46, 8'h19, 8'h0, 8'hd, 8'h31, 8'h65, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h5d, 8'h2b, 8'h32, 8'h7b, 8'h7e, 8'h27, 8'h0, 8'h37, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h8f, 8'h78, 8'h4a, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3b, 8'h53, 8'h77, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h45, 8'h0, 8'h4c, 8'h88, 8'h9a, 8'h99, 8'h96, 8'h92, 8'h87, 8'h73, 8'h50, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7c, 8'h7, 8'h0, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h63, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h1d, 8'h8, 8'h77, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h61, 8'h7, 8'h0, 8'h60, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h37, 8'h0, 8'h0, 8'h4a, 8'h8b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h3b, 8'h0, 8'h0, 8'h58, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h44, 8'h0, 8'h23, 8'h74, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h68, 8'h0, 8'h0, 8'h27, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h88, 8'h30, 8'h0, 8'h0, 8'h1, 8'h45, 8'h74, 8'h81, 8'h3c, 8'h0, 8'h4d, 8'h88, 8'h9a, 8'h90, 8'h5c, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h68, 8'h3, 8'h0, 8'h50, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6d, 8'h16, 8'h11, 8'h85, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7c, 8'h31, 8'h0, 8'h46, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h4d, 8'h9, 8'h1b, 8'h5a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h97, 8'h8b, 8'h68, 8'h24, 8'ha, 8'h0, 8'h17, 8'h62, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h86, 8'h87, 8'h99, 8'h7d, 8'h14, 8'hb, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h91, 8'h87, 8'h6f, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h62, 8'h7c, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h42, 8'h0, 8'h50, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h8d, 8'h6c, 8'h26, 8'h0, 8'h0, 8'h0, 8'h9, 8'h70, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h75, 8'h0, 8'h12, 8'h64, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h6d, 8'h45, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h76, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7b, 8'h29, 8'h0, 8'h59, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h41, 8'h0, 8'h0, 8'h2d, 8'h70, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h40, 8'h0, 8'h0, 8'h54, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h42, 8'h0, 8'h16, 8'h6e, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h61, 8'h0, 8'h0, 8'h32, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h40, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h4b, 8'h20, 8'h0, 8'h5c, 8'h8c, 8'h9b, 8'h95, 8'h65, 8'h0, 8'h0, 8'h36, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h69, 8'h5, 8'h0, 8'h51, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h54, 8'h12, 8'h27, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h4b, 8'h0, 8'h16, 8'h6a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h4c, 8'h0, 8'hd, 8'h5b, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h89, 8'h69, 8'h1e, 8'h0, 8'h5, 8'h6a, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7b, 8'hc, 8'h11, 8'h6f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h8c, 8'h7a, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h77, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h3b, 8'h0, 8'h5e, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7c, 8'h29, 8'h0, 8'h0, 8'h0, 8'h7, 8'h78, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h69, 8'h0, 8'h3a, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h74, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7c, 8'h2d, 8'h0, 8'h59, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h69, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h85, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8e, 8'h3e, 8'h0, 8'h0, 8'h51, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h3c, 8'h0, 8'h5, 8'h65, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h66, 8'h0, 8'h0, 8'h29, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h7b, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7a, 8'h99, 8'h9a, 8'h98, 8'h6a, 8'h0, 8'h0, 8'h31, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h80, 8'h39, 8'h0, 8'h48, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h70, 8'h49, 8'h5a, 8'h9b, 8'h9b, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h5f, 8'hb, 8'h0, 8'h65, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h49, 8'h0, 8'h0, 8'h6a, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h7c, 8'h2c, 8'h0, 8'h0, 8'h69, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6d, 8'h7, 8'h22, 8'h85, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h88, 8'h6e, 8'h54, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h71, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h80, 8'h2f, 8'h0, 8'h64, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7a, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h5e, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7c, 8'h2d, 8'h0, 8'h48, 8'h98, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h8b, 8'h85, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h7b, 8'h4d, 8'h15, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h4c, 8'h59, 8'h5a, 8'h59, 8'h63, 8'h7a, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h32, 8'h0, 8'h56, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h56, 8'h31, 8'h41, 8'h7b, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h41, 8'h0, 8'h0, 8'h47, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h39, 8'h0, 8'h0, 8'h62, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7b, 8'h1f, 8'h0, 8'h0, 8'h4f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h7c, 8'h64, 8'h58, 8'h47, 8'h22, 8'hd, 8'h20, 8'h5f, 8'h91, 8'h9b, 8'h9b, 8'h99, 8'h6b, 8'h0, 8'h0, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h63, 8'h0, 8'h25, 8'h77, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h85, 8'h89, 8'h9a, 8'h87, 8'h3c, 8'h41, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h61, 8'h18, 8'h0, 8'h32, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h61, 8'h16, 8'h2, 8'h5a, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h79, 8'h32, 8'h0, 8'h8, 8'h5d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h56, 8'h0, 8'h2c, 8'h94, 8'h93, 8'h6b, 8'h39, 8'h26, 8'h4d, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h92, 8'h7e, 8'h50, 8'h23, 8'h0, 8'h0, 8'h0, 8'hb, 8'h4b, 8'h80, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6e, 8'h16, 8'h0, 8'h6a, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h5f, 8'h34, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h55, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h63, 8'h0, 8'h0, 8'h56, 8'h90, 8'h76, 8'h44, 8'h2e, 8'h2b, 8'h26, 8'h2a, 8'h62, 8'h8d, 8'h9a, 8'h99, 8'h82, 8'h36, 8'h1, 8'h0, 8'h0, 8'h1b, 8'h34, 8'h5d, 8'h7d, 8'h90, 8'h95, 8'h95, 8'h94, 8'h96, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h35, 8'h0, 8'h4a, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h8d, 8'h85, 8'h7d, 8'h79, 8'h74, 8'h6f, 8'h6b, 8'h6b, 8'h67, 8'h65, 8'h64, 8'h65, 8'h64, 8'h64, 8'h63, 8'h62, 8'h60, 8'h61, 8'h64, 8'h65, 8'h65, 8'h65, 8'h64, 8'h5f, 8'h52, 8'h43, 8'h47, 8'h60, 8'h64, 8'h62, 8'h64, 8'h64, 8'h62, 8'h61, 8'h57, 8'h24, 8'h0, 8'h0, 8'hf, 8'h4c, 8'h66, 8'h65, 8'h6a, 8'h6c, 8'h70, 8'h73, 8'h78, 8'h81, 8'h86, 8'h7a, 8'h33, 8'h0, 8'h0, 8'h5d, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h55, 8'h0, 8'h0, 8'h28, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h97, 8'h94, 8'h8d, 8'h74, 8'h65, 8'h71, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h98, 8'h6e, 8'h0, 8'h0, 8'h2a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h78, 8'h4, 8'h3, 8'h4f, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h99, 8'h9b, 8'h80, 8'h16, 8'h0, 8'h3a, 8'h90, 8'h99, 8'h9b, 8'h97, 8'h7a, 8'h3e, 8'h1d, 8'h0, 8'h0, 8'h1d, 8'h73, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h7e, 8'h2a, 8'h9, 8'h39, 8'h8e, 8'h97, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h79, 8'h2e, 8'h0, 8'hb, 8'h57, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h42, 8'h0, 8'h2f, 8'h88, 8'h5c, 8'h16, 8'h0, 8'h0, 8'h2d, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h91, 8'h7e, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h5e, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5a, 8'h0, 8'h0, 8'h6a, 8'h7c, 8'h76, 8'h87, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h8e, 8'h7e, 8'h51, 8'hf, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h61, 8'h86, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h54, 8'h0, 8'h3, 8'h36, 8'h46, 8'h23, 8'h0, 8'h1, 8'h11, 8'h0, 8'h0, 8'h15, 8'h74, 8'h9b, 8'h99, 8'h7b, 8'h1b, 8'h0, 8'h0, 8'h49, 8'h7c, 8'h8c, 8'h95, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h3d, 8'h0, 8'h1f, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h8c, 8'h84, 8'h7e, 8'h79, 8'h76, 8'h75, 8'h76, 8'h76, 8'h76, 8'h77, 8'h78, 8'h78, 8'h75, 8'h73, 8'h6d, 8'h68, 8'h6a, 8'h68, 8'h65, 8'h63, 8'h62, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h5c, 8'h5a, 8'h58, 8'h57, 8'h58, 8'h5b, 8'h5c, 8'h5d, 8'h5d, 8'h5c, 8'h5a, 8'h5a, 8'h59, 8'h5a, 8'h5e, 8'h5b, 8'h5b, 8'h5b, 8'h5c, 8'h58, 8'h57, 8'h54, 8'h3d, 8'hd, 8'h0, 8'h1c, 8'h48, 8'h5d, 8'h5d, 8'h61, 8'h64, 8'h65, 8'h65, 8'h66, 8'h6d, 8'h6e, 8'h63, 8'h25, 8'h0, 8'h0, 8'h3f, 8'h76, 8'h74, 8'h75, 8'h77, 8'h79, 8'h7c, 8'h80, 8'h88, 8'h8e, 8'h94, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7d, 8'h14, 8'h0, 8'h0, 8'h49, 8'h5f, 8'h85, 8'h94, 8'h96, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h95, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h7c, 8'h8, 8'h0, 8'h3c, 8'h94, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h88, 8'h35, 8'h0, 8'h25, 8'h80, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h35, 8'h0, 8'h0, 8'h4d, 8'h8b, 8'h9a, 8'h93, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h43, 8'h6, 8'h24, 8'h72, 8'h99, 8'h9b, 8'h9a, 8'h98, 8'h86, 8'h5c, 8'h53, 8'h5b, 8'h79, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7a, 8'h2c, 8'h0, 8'h7, 8'h54, 8'h7c, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h3a, 8'h0, 8'h1c, 8'h4f, 8'h0, 8'h0, 8'h0, 8'he, 8'h62, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h85, 8'h6f, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h4a, 8'h0, 8'h0, 8'h49, 8'h37, 8'h29, 8'h5a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h7f, 8'h52, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h47, 8'h78, 8'h8d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h50, 8'h0, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4b, 8'h70, 8'h44, 8'h0, 8'h0, 8'h4d, 8'h8f, 8'h99, 8'h88, 8'h40, 8'h0, 8'h8, 8'h64, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h4c, 8'h0, 8'h0, 8'h51, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h94, 8'h90, 8'h8c, 8'h8a, 8'h8a, 8'h89, 8'h89, 8'h8a, 8'h88, 8'h80, 8'h71, 8'h64, 8'h59, 8'h51, 8'h4b, 8'h48, 8'h49, 8'h49, 8'h49, 8'h4b, 8'h4f, 8'h53, 8'h58, 8'h61, 8'h6a, 8'h73, 8'h81, 8'h89, 8'h8e, 8'h91, 8'h93, 8'h92, 8'h93, 8'h93, 8'h94, 8'h92, 8'h93, 8'h92, 8'h92, 8'h92, 8'h92, 8'h93, 8'h93, 8'h93, 8'h92, 8'h93, 8'h92, 8'h93, 8'h93, 8'h93, 8'h92, 8'h93, 8'h93, 8'h93, 8'h93, 8'h92, 8'h91, 8'h92, 8'h8f, 8'h7a, 8'h59, 8'h78, 8'h8e, 8'h92, 8'h93, 8'h92, 8'h92, 8'h8d, 8'h85, 8'h79, 8'h74, 8'h69, 8'h5a, 8'h2a, 8'h0, 8'h0, 8'h2b, 8'h4b, 8'h46, 8'h47, 8'h4c, 8'h50, 8'h55, 8'h5c, 8'h6b, 8'h77, 8'h7f, 8'h85, 8'h8a, 8'h8b, 8'h8a, 8'h8a, 8'h8b, 8'h8d, 8'h90, 8'h94, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h64, 8'hf, 8'h0, 8'h0, 8'h0, 8'h47, 8'h6a, 8'h6c, 8'h70, 8'h75, 8'h79, 8'h81, 8'h89, 8'h90, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h5d, 8'h36, 8'h40, 8'h68, 8'h72, 8'h7e, 8'h8f, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7a, 8'h23, 8'h9, 8'h47, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h8a, 8'h85, 8'h81, 8'h85, 8'h8f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h1a, 8'h0, 8'h0, 8'h66, 8'h91, 8'h95, 8'h6b, 8'h15, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8b, 8'h55, 8'h0, 8'he, 8'h5a, 8'h97, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h30, 8'h0, 8'h0, 8'h35, 8'h6e, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h6e, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h79, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h1, 8'h45, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h7d, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h53, 8'h0, 8'h0, 8'h0, 8'hb, 8'h66, 8'h82, 8'h91, 8'h95, 8'h7c, 8'h2c, 8'h0, 8'h0, 8'h5b, 8'h9b, 8'h99, 8'h73, 8'h0, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h4e, 8'h0, 8'h0, 8'h49, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8b, 8'h76, 8'h5d, 8'h48, 8'h41, 8'h3e, 8'h3c, 8'h3b, 8'h43, 8'h4a, 8'h55, 8'h64, 8'h78, 8'h85, 8'h8b, 8'h8c, 8'h8d, 8'h8d, 8'h8e, 8'h8e, 8'h8e, 8'h8e, 8'h8f, 8'h91, 8'h91, 8'h93, 8'h95, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h94, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h95, 8'h95, 8'h91, 8'h86, 8'h74, 8'h7c, 8'h89, 8'h8e, 8'h8d, 8'h8d, 8'h8e, 8'h8e, 8'h8b, 8'h85, 8'h76, 8'h66, 8'h53, 8'h45, 8'h42, 8'h40, 8'h3f, 8'h3f, 8'h43, 8'h4d, 8'h5e, 8'h76, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h7a, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h3b, 8'h60, 8'h82, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7e, 8'h17, 8'h0, 8'h0, 8'h0, 8'h4, 8'h5a, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h75, 8'h35, 8'hf, 8'h52, 8'h8a, 8'h9a, 8'h9b, 8'h95, 8'h7f, 8'h45, 8'h1e, 8'h11, 8'h27, 8'h5e, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h66, 8'h10, 8'h0, 8'h20, 8'h75, 8'h9b, 8'h94, 8'h87, 8'h80, 8'h6f, 8'h29, 8'h0, 8'h51, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h4e, 8'h0, 8'h0, 8'h58, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h8e, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h41, 8'h0, 8'h0, 8'h4, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7e, 8'h13, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h48, 8'h2e, 8'h34, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h85, 8'h4c, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h68, 8'h74, 8'h6b, 8'h82, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h92, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h69, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4, 8'h2a, 8'h68, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h75, 8'h20, 8'h0, 8'h1c, 8'h6a, 8'h91, 8'h99, 8'h9b, 8'h9a, 8'h8f, 8'h59, 8'h0, 8'h0, 8'h49, 8'h9b, 8'h9a, 8'h85, 8'h25, 8'h0, 8'h12, 8'h95, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h4f, 8'h0, 8'h0, 8'h46, 8'h95, 8'h87, 8'h73, 8'h63, 8'h5a, 8'h55, 8'h54, 8'h56, 8'h5b, 8'h63, 8'h6d, 8'h75, 8'h77, 8'h79, 8'h78, 8'h78, 8'h77, 8'h7a, 8'h7d, 8'h82, 8'h88, 8'h91, 8'h97, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h90, 8'h89, 8'h81, 8'h7b, 8'h7a, 8'h78, 8'h79, 8'h79, 8'h79, 8'h79, 8'h71, 8'h69, 8'h62, 8'h5a, 8'h53, 8'h55, 8'h56, 8'h59, 8'h63, 8'h74, 8'h8b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h82, 8'h64, 8'h59, 8'h57, 8'h55, 8'h54, 8'h50, 8'h3a, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h1b, 8'h3f, 8'h62, 8'h7c, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h6a, 8'h47, 8'h27, 8'h0, 8'h0, 8'h0, 8'h3, 8'h33, 8'h83, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h80, 8'h61, 8'h4e, 8'h71, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h7d, 8'h6a, 8'h81, 8'h94, 8'h92, 8'h5b, 8'hc, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h40, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h40, 8'h0, 8'h0, 8'h5c, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h65, 8'h1e, 8'hd, 8'h79, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h46, 8'h0, 8'h0, 8'h54, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h77, 8'h2b, 8'h7, 8'h5c, 8'h52, 8'h2c, 8'h0, 8'h0, 8'h28, 8'h80, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h53, 8'h1c, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h73, 8'h0, 8'h0, 8'h0, 8'h2, 8'h44, 8'h70, 8'h34, 8'h0, 8'ha, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h85, 8'h57, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h52, 8'h80, 8'h94, 8'h97, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h76, 8'hd, 8'h0, 8'h0, 8'hd, 8'h4, 8'h0, 8'h7, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h96, 8'h86, 8'h5a, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9, 8'h5b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h6c, 8'h45, 8'h6a, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h79, 8'h1e, 8'h0, 8'h36, 8'h8e, 8'h9b, 8'h91, 8'h58, 8'h1, 8'h0, 8'h6d, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h89, 8'h75, 8'h30, 8'h0, 8'h0, 8'h26, 8'h69, 8'h6a, 8'h6b, 8'h6b, 8'h6b, 8'h68, 8'h68, 8'h6a, 8'h6f, 8'h77, 8'h82, 8'h8e, 8'h94, 8'h97, 8'h98, 8'h99, 8'h98, 8'h98, 8'h98, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h98, 8'h98, 8'h98, 8'h99, 8'h98, 8'h98, 8'h95, 8'h8c, 8'h7f, 8'h75, 8'h6d, 8'h67, 8'h69, 8'h69, 8'h6b, 8'h6c, 8'h68, 8'h69, 8'h69, 8'h68, 8'h66, 8'h69, 8'h6f, 8'h7b, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h95, 8'h96, 8'h95, 8'h94, 8'h91, 8'h83, 8'h5c, 8'h3b, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h26, 8'h33, 8'h43, 8'h61, 8'h80, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h8c, 8'h77, 8'h4b, 8'h20, 8'h0, 8'h0, 8'h0, 8'h20, 8'h5b, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h59, 8'h26, 8'h14, 8'h0, 8'h0, 8'h49, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h96, 8'h99, 8'h95, 8'h70, 8'h1c, 8'h0, 8'h0, 8'hd, 8'h28, 8'h2c, 8'h2c, 8'h2f, 8'h5c, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h73, 8'h22, 8'h0, 8'h3b, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h47, 8'h0, 8'h3f, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h45, 8'h1, 8'h0, 8'h4a, 8'h89, 8'h9a, 8'h9a, 8'h9b, 8'h98, 8'h82, 8'h3f, 8'h13, 8'h34, 8'h93, 8'h91, 8'h78, 8'h43, 8'h0, 8'h0, 8'h39, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8d, 8'h68, 8'h28, 8'h0, 8'h0, 8'h50, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h78, 8'hb, 8'h0, 8'h1b, 8'h5b, 8'h91, 8'h7f, 8'h11, 8'h0, 8'h9, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h91, 8'h69, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h51, 8'h8a, 8'h93, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h68, 8'h6, 8'h0, 8'h19, 8'h63, 8'h36, 8'h0, 8'h8, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h7a, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h91, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8f, 8'h58, 8'h0, 8'hd, 8'h63, 8'h9b, 8'h97, 8'h79, 8'h16, 8'h0, 8'h2c, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h8b, 8'h82, 8'h7b, 8'h79, 8'h78, 8'h77, 8'h70, 8'h60, 8'h27, 8'h0, 8'h0, 8'h1e, 8'h60, 8'h6d, 8'h7f, 8'h8c, 8'h93, 8'h95, 8'h95, 8'h95, 8'h96, 8'h97, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h96, 8'h95, 8'h95, 8'h96, 8'h95, 8'h94, 8'h8c, 8'h7a, 8'h69, 8'h5f, 8'h5a, 8'h59, 8'h5c, 8'h60, 8'h67, 8'h71, 8'h7c, 8'h79, 8'h78, 8'h7b, 8'h81, 8'h8c, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h71, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h2, 8'h0, 8'h0, 8'he, 8'h31, 8'h4d, 8'h5a, 8'h66, 8'h7f, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h91, 8'h7b, 8'h38, 8'h0, 8'h0, 8'h0, 8'h3, 8'h46, 8'h7d, 8'h9b, 8'h9a, 8'h7f, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h5, 8'h54, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h8d, 8'h41, 8'h0, 8'h0, 8'h1d, 8'h6b, 8'h8a, 8'h8d, 8'h8d, 8'h88, 8'h8e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h62, 8'h0, 8'h17, 8'h6a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6c, 8'h17, 8'h10, 8'h61, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8c, 8'h51, 8'h0, 8'h0, 8'h40, 8'h91, 8'h99, 8'h9a, 8'h9b, 8'h98, 8'h87, 8'h47, 8'h12, 8'h24, 8'h6a, 8'h99, 8'h9b, 8'h97, 8'h84, 8'h48, 8'h0, 8'h0, 8'h51, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h72, 8'h2c, 8'h0, 8'h0, 8'h53, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7f, 8'h81, 8'h8a, 8'h94, 8'h9b, 8'h7e, 8'h2, 8'h0, 8'h6, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h89, 8'h61, 8'h9, 8'h0, 8'h0, 8'h0, 8'h6, 8'h60, 8'h87, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h70, 8'h24, 8'h18, 8'h85, 8'h88, 8'h47, 8'h0, 8'h6, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h7b, 8'h46, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h79, 8'h2, 8'h0, 8'h23, 8'h95, 8'h9a, 8'h86, 8'h26, 8'h0, 8'h0, 8'h7c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h90, 8'h8d, 8'h8d, 8'h8c, 8'h84, 8'h6c, 8'h59, 8'h4c, 8'h46, 8'h46, 8'h51, 8'h63, 8'h72, 8'h4e, 8'h0, 8'h0, 8'h51, 8'h93, 8'h95, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h94, 8'h92, 8'h92, 8'h92, 8'h92, 8'h8e, 8'h7a, 8'h63, 8'h51, 8'h49, 8'h46, 8'h4b, 8'h5b, 8'h6f, 8'h85, 8'h8b, 8'h8d, 8'h8d, 8'h90, 8'h96, 8'h8e, 8'h52, 8'h0, 8'h0, 8'h39, 8'h67, 8'h53, 8'h8, 8'h0, 8'h58, 8'h7c, 8'h69, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h64, 8'h79, 8'h7e, 8'h81, 8'h8d, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8d, 8'h7a, 8'h40, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h8f, 8'h98, 8'h7e, 8'h24, 8'h0, 8'h6, 8'h3e, 8'h70, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h82, 8'h14, 8'h0, 8'h0, 8'h7c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h6e, 8'h0, 8'h0, 8'h56, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h66, 8'ha, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h90, 8'h63, 8'h0, 8'h0, 8'h3f, 8'h8c, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h89, 8'h52, 8'h0, 8'h1a, 8'h62, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h73, 8'h17, 8'h0, 8'h2d, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h76, 8'h30, 8'h0, 8'h0, 8'h52, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h7e, 8'h0, 8'h0, 8'h8, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h80, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h50, 8'h7e, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h87, 8'h84, 8'h9a, 8'h91, 8'h54, 8'h5, 8'h4, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h65, 8'h8, 8'h0, 8'h0, 8'h0, 8'h16, 8'h61, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8b, 8'h41, 8'h0, 8'h5, 8'h7a, 8'h96, 8'h8e, 8'h52, 8'h0, 8'h0, 8'h65, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h93, 8'h7b, 8'h59, 8'h47, 8'h44, 8'h45, 8'h52, 8'h67, 8'h7e, 8'h89, 8'h8a, 8'h89, 8'h8d, 8'h90, 8'h94, 8'h8b, 8'h72, 8'h76, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h91, 8'h8c, 8'h8a, 8'h8a, 8'h89, 8'h7a, 8'h64, 8'h4f, 8'h41, 8'h3f, 8'h45, 8'h57, 8'h78, 8'h85, 8'h4b, 8'h0, 8'h0, 8'h44, 8'h71, 8'h38, 8'h0, 8'h0, 8'h74, 8'h97, 8'h96, 8'h8b, 8'h7d, 8'h79, 8'h6b, 8'h4a, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3f, 8'h74, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8c, 8'h60, 8'h4, 8'h0, 8'h0, 8'h4d, 8'h92, 8'h97, 8'h86, 8'h7c, 8'h81, 8'h8c, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h80, 8'h8, 8'h0, 8'h0, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h69, 8'h0, 8'h1a, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h76, 8'he, 8'h53, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6c, 8'h18, 8'h0, 8'h3e, 8'h84, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h58, 8'h0, 8'h3, 8'h5a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6e, 8'hb, 8'h0, 8'h30, 8'h84, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h95, 8'h7d, 8'h3e, 8'h0, 8'h0, 8'h4c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h0, 8'h0, 8'hf, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h61, 8'h88, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h91, 8'h5f, 8'hd, 8'h3, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h77, 8'h56, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h41, 8'h6e, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h6e, 8'ha, 8'h0, 8'h35, 8'h8c, 8'h98, 8'h7a, 8'h25, 8'h0, 8'h17, 8'h72, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h74, 8'h5f, 8'h58, 8'h59, 8'h5f, 8'h6a, 8'h70, 8'h74, 8'h78, 8'h78, 8'h7c, 8'h88, 8'h94, 8'h99, 8'h9a, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h95, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h99, 8'h92, 8'h87, 8'h7d, 8'h76, 8'h74, 8'h75, 8'h71, 8'h63, 8'h57, 8'h38, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h94, 8'h86, 8'h6e, 8'h56, 8'h4e, 8'h3f, 8'h27, 8'h1, 8'h0, 8'h0, 8'h0, 8'h8, 8'h17, 8'h2e, 8'h55, 8'h81, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h59, 8'h0, 8'h0, 8'h11, 8'h8c, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h7, 8'h0, 8'h0, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h67, 8'he, 8'h0, 8'h46, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h77, 8'h7, 8'h50, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7b, 8'h35, 8'h0, 8'h1e, 8'h72, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h64, 8'h13, 8'h0, 8'h4d, 8'h88, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h73, 8'h29, 8'h0, 8'h1a, 8'h64, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h7c, 8'h35, 8'h0, 8'h0, 8'h43, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h0, 8'h0, 8'h1a, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h63, 8'ha, 8'h0, 8'h0, 8'h34, 8'h72, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5d, 8'hb, 8'h2, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h78, 8'h32, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h4e, 8'h88, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h22, 8'h0, 8'h3, 8'h82, 8'h98, 8'h8e, 8'h46, 8'h0, 8'h0, 8'h43, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h7c, 8'h6e, 8'h6b, 8'h6c, 8'h6c, 8'h69, 8'h6a, 8'h66, 8'h67, 8'h6e, 8'h7c, 8'h8d, 8'h95, 8'h97, 8'h98, 8'h98, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h97, 8'h97, 8'h95, 8'h8d, 8'h79, 8'h6d, 8'h61, 8'h46, 8'h19, 8'h0, 8'h0, 8'h0, 8'ha, 8'h4f, 8'h78, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h97, 8'h95, 8'h91, 8'h8a, 8'h76, 8'h57, 8'h34, 8'h26, 8'h16, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h48, 8'h72, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7d, 8'h8, 8'h0, 8'h0, 8'h8a, 8'h9b, 8'h9a, 8'h95, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h80, 8'h5, 8'h0, 8'h0, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h7f, 8'h51, 8'h11, 8'h0, 8'h25, 8'h75, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h75, 8'h7, 8'h50, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h98, 8'h80, 8'h41, 8'h1, 8'h1, 8'h60, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3b, 8'h0, 8'h1b, 8'h7d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h71, 8'h31, 8'h0, 8'hf, 8'h5b, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7a, 8'h35, 8'h0, 8'h0, 8'h42, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h76, 8'h0, 8'h0, 8'h29, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h61, 8'h2b, 8'h0, 8'h0, 8'h43, 8'h81, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h52, 8'h3, 8'h4, 8'h91, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h7b, 8'h70, 8'h85, 8'h9a, 8'h9b, 8'h96, 8'h6c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h38, 8'h72, 8'h94, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h4a, 8'h0, 8'h0, 8'h62, 8'h8f, 8'h94, 8'h66, 8'h7, 8'h0, 8'h8, 8'h61, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h8a, 8'h80, 8'h7e, 8'h7d, 8'h75, 8'h64, 8'h5b, 8'h57, 8'h5b, 8'h68, 8'h7c, 8'h90, 8'h94, 8'h95, 8'h96, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h97, 8'h95, 8'h94, 8'h91, 8'h81, 8'h5a, 8'h33, 8'h30, 8'h45, 8'h58, 8'h66, 8'h76, 8'h7c, 8'h7e, 8'h81, 8'h8b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h92, 8'h8f, 8'h89, 8'h75, 8'h4c, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h4e, 8'h62, 8'h7b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h78, 8'h5, 8'h0, 8'h0, 8'h8b, 8'h99, 8'h8c, 8'h6c, 8'h48, 8'h60, 8'h83, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7f, 8'h8, 8'h0, 8'h0, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h72, 8'h5f, 8'h59, 8'h59, 8'h53, 8'h34, 8'h0, 8'h0, 8'h15, 8'h70, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h6b, 8'h7, 8'h51, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h4b, 8'h6, 8'h0, 8'h46, 8'h8b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h85, 8'h24, 8'h0, 8'h3b, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h77, 8'h35, 8'h1, 8'hb, 8'h5a, 8'h8b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7c, 8'h37, 8'h0, 8'h0, 8'h47, 8'h81, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6e, 8'h0, 8'h0, 8'h3c, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h86, 8'h33, 8'h0, 8'h4, 8'h5a, 8'h8f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h47, 8'h0, 8'h8, 8'h91, 8'h9a, 8'h91, 8'h83, 8'h63, 8'h2b, 8'h9, 8'h47, 8'h8d, 8'h9b, 8'h9a, 8'h7d, 8'he, 8'h0, 8'h0, 8'h53, 8'h86, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h2b, 8'h0, 8'h21, 8'h78, 8'h9a, 8'h8f, 8'h59, 8'h0, 8'h0, 8'h2d, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h93, 8'h90, 8'h8d, 8'h82, 8'h66, 8'h4d, 8'h47, 8'h4d, 8'h59, 8'h72, 8'h8f, 8'h91, 8'h92, 8'h94, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h90, 8'h8e, 8'h91, 8'h8b, 8'h73, 8'h58, 8'h4a, 8'h49, 8'h51, 8'h69, 8'h83, 8'h91, 8'h90, 8'h92, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h92, 8'h8b, 8'h82, 8'h64, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h6d, 8'h87, 8'h8b, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h60, 8'h0, 8'h0, 8'h1d, 8'h8d, 8'h96, 8'h76, 8'h24, 8'h0, 8'h0, 8'h49, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h80, 8'ha, 8'h0, 8'h0, 8'h8b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h23, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h83, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h4f, 8'h5, 8'h53, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h91, 8'h62, 8'h0, 8'h0, 8'h3c, 8'h91, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h29, 8'h0, 8'hd, 8'h74, 8'h94, 8'h9a, 8'h99, 8'h85, 8'h3b, 8'h0, 8'hb, 8'h5a, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h40, 8'h0, 8'h0, 8'h43, 8'h87, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h66, 8'h0, 8'h0, 8'h4e, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h66, 8'h0, 8'h0, 8'h17, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8c, 8'h46, 8'h0, 8'h6, 8'h93, 8'h90, 8'h59, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h9b, 8'h9a, 8'h8f, 8'h55, 8'h0, 8'h0, 8'h19, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h3b, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h99, 8'h80, 8'h23, 8'h0, 8'h0, 8'h4e, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h7f, 8'h5b, 8'h4b, 8'h49, 8'h51, 8'h66, 8'h80, 8'h86, 8'h88, 8'h8c, 8'h92, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h8c, 8'h87, 8'h87, 8'h82, 8'h64, 8'h50, 8'h45, 8'h4b, 8'h60, 8'h82, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h7f, 8'h66, 8'h44, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h55, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7e, 8'hb, 8'h0, 8'h0, 8'h69, 8'h96, 8'h99, 8'h8a, 8'h44, 8'h0, 8'h0, 8'h15, 8'h6c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hf, 8'h0, 8'h0, 8'h8c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h58, 8'h84, 8'h98, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6e, 8'h15, 8'h8, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h6b, 8'h0, 8'h0, 8'h3b, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h93, 8'h60, 8'hc, 8'h0, 8'hc, 8'h6c, 8'h9a, 8'h8a, 8'h55, 8'h0, 8'hc, 8'h53, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h4d, 8'h0, 8'h0, 8'h38, 8'h8f, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h58, 8'h0, 8'h0, 8'h5f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h28, 8'h0, 8'h0, 8'h2b, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h50, 8'h1, 8'h5, 8'h83, 8'h4a, 8'h3, 8'h0, 8'h0, 8'h21, 8'h0, 8'h0, 8'h18, 8'h87, 8'h98, 8'h99, 8'h7d, 8'h26, 8'h0, 8'h0, 8'h5e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h66, 8'h9, 8'h0, 8'h3f, 8'h88, 8'h9b, 8'h92, 8'h69, 8'h12, 8'h0, 8'h27, 8'h80, 8'h64, 8'h5b, 8'h5c, 8'h64, 8'h70, 8'h74, 8'h73, 8'h7b, 8'h87, 8'h96, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h86, 8'h7b, 8'h72, 8'h71, 8'h6e, 8'h64, 8'h5d, 8'h5c, 8'h67, 8'h81, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h85, 8'h68, 8'h48, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h35, 8'h78, 8'h96, 8'h99, 8'h91, 8'h60, 8'h0, 8'h0, 8'h1d, 8'h8e, 8'h9a, 8'h9b, 8'h96, 8'h7d, 8'h54, 8'h4a, 8'h63, 8'h85, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h1e, 8'h0, 8'h0, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h5a, 8'h41, 8'h44, 8'h52, 8'h71, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h58, 8'h0, 8'h3b, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h69, 8'h17, 8'h0, 8'h35, 8'h79, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h5e, 8'h18, 8'h0, 8'h10, 8'h53, 8'h5d, 8'h0, 8'h0, 8'h3e, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h75, 8'h50, 8'h4e, 8'h7f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h42, 8'h0, 8'h0, 8'h33, 8'h85, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h35, 8'h0, 8'ha, 8'h72, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h90, 8'h94, 8'h97, 8'h8a, 8'h64, 8'h49, 8'h8d, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h61, 8'h8, 8'h0, 8'h0, 8'h5d, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5c, 8'h9, 8'h0, 8'h47, 8'h1, 8'h0, 8'h0, 8'h4a, 8'h72, 8'h2c, 8'h0, 8'h0, 8'h46, 8'h92, 8'h9a, 8'h8f, 8'h50, 8'h0, 8'h0, 8'h24, 8'h75, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h46, 8'h0, 8'h6, 8'h5d, 8'h98, 8'h96, 8'h74, 8'h37, 8'h13, 8'h2a, 8'h67, 8'h66, 8'h64, 8'h66, 8'h77, 8'h8d, 8'h95, 8'h98, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h97, 8'h98, 8'h94, 8'h89, 8'h74, 8'h68, 8'h64, 8'h67, 8'h6a, 8'h6d, 8'h6e, 8'h73, 8'h84, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h8e, 8'h6e, 8'h3f, 8'h1a, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h40, 8'h66, 8'h6c, 8'h15, 8'h0, 8'h0, 8'h50, 8'h98, 8'h87, 8'h5f, 8'h75, 8'h95, 8'h94, 8'h94, 8'h95, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h40, 8'h0, 8'h0, 8'h5b, 8'h8d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h95, 8'h92, 8'h92, 8'h93, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h7a, 8'h30, 8'h0, 8'h64, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6b, 8'h24, 8'h0, 8'h18, 8'h6f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8e, 8'h65, 8'h15, 8'h0, 8'h0, 8'h6, 8'h0, 8'h1, 8'h60, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h84, 8'h48, 8'h1c, 8'h0, 8'h0, 8'h2b, 8'h66, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h84, 8'h41, 8'h0, 8'h0, 8'h33, 8'h7a, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7f, 8'ha, 8'h0, 8'h17, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h88, 8'h6f, 8'h55, 8'h4e, 8'h64, 8'h82, 8'h77, 8'h30, 8'h0, 8'h65, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h41, 8'h0, 8'h0, 8'h21, 8'h73, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h5b, 8'h1, 8'h0, 8'h0, 8'h0, 8'h6, 8'h54, 8'h92, 8'h97, 8'h71, 8'h4, 8'h0, 8'h5, 8'h85, 8'h9b, 8'h96, 8'h75, 8'h26, 8'h0, 8'h0, 8'h43, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h6f, 8'h0, 8'h0, 8'h2f, 8'h7d, 8'h79, 8'h67, 8'h53, 8'h48, 8'h52, 8'h6f, 8'h8b, 8'h93, 8'h95, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h94, 8'h94, 8'h8a, 8'h6e, 8'h5b, 8'h54, 8'h5a, 8'h68, 8'h7c, 8'h82, 8'h86, 8'h8f, 8'h9a, 8'h9b, 8'h99, 8'h95, 8'h88, 8'h6b, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h20, 8'h0, 8'h0, 8'h2e, 8'h84, 8'h97, 8'h75, 8'h17, 8'h37, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6a, 8'h10, 8'h0, 8'h1a, 8'h77, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h7c, 8'h74, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h89, 8'h4c, 8'h9, 8'h17, 8'h7b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h79, 8'h2d, 8'h0, 8'h4, 8'h63, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h92, 8'h67, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h34, 8'h78, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h66, 8'h91, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h49, 8'h0, 8'h0, 8'h37, 8'h79, 8'h96, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h76, 8'h0, 8'h0, 8'h24, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h82, 8'h4e, 8'h3, 8'h0, 8'h0, 8'h7, 8'h60, 8'h7f, 8'h3b, 8'h0, 8'h21, 8'h75, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h81, 8'h33, 8'h0, 8'h0, 8'h47, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8a, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h94, 8'h9b, 8'h9b, 8'h82, 8'h16, 8'h0, 8'h0, 8'h70, 8'h93, 8'h99, 8'h94, 8'h63, 8'h0, 8'h0, 8'h1a, 8'h7a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h95, 8'h89, 8'h5c, 8'h14, 8'h1b, 8'h42, 8'h4c, 8'h6c, 8'h87, 8'h92, 8'h91, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h95, 8'h92, 8'h8f, 8'h82, 8'h67, 8'h4b, 8'h48, 8'h54, 8'h72, 8'h92, 8'h93, 8'h95, 8'h94, 8'h78, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h99, 8'h9b, 8'h7b, 8'ha, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h2e, 8'h0, 8'h0, 8'h58, 8'h90, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h79, 8'h2d, 8'h17, 8'h8a, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h8c, 8'h65, 8'h1c, 8'h0, 8'h5b, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h44, 8'h0, 8'h0, 8'h53, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h82, 8'h72, 8'h71, 8'h85, 8'h8e, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h66, 8'h13, 8'h0, 8'h0, 8'h43, 8'h57, 8'h3, 8'h0, 8'h22, 8'h6f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h51, 8'h0, 8'h0, 8'h3b, 8'h86, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h73, 8'h0, 8'h0, 8'h29, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6b, 8'h0, 8'h0, 8'h0, 8'hd, 8'h65, 8'h75, 8'h8a, 8'h8f, 8'h57, 8'h0, 8'h0, 8'h5a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5b, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h4, 8'h0, 8'h0, 8'he, 8'h60, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h52, 8'h0, 8'h0, 8'h10, 8'h75, 8'h9b, 8'h9a, 8'h89, 8'h41, 8'h0, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h78, 8'h58, 8'h4a, 8'h49, 8'h54, 8'h6e, 8'h84, 8'h85, 8'h90, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8f, 8'h86, 8'h83, 8'h78, 8'h64, 8'h4e, 8'h4d, 8'h5f, 8'h75, 8'h4b, 8'h0, 8'h0, 8'h43, 8'h68, 8'h2e, 8'h0, 8'h0, 8'h2a, 8'h18, 8'h0, 8'h0, 8'h4b, 8'h89, 8'h9b, 8'h9b, 8'h89, 8'h39, 8'h0, 8'h27, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h64, 8'ha, 8'h0, 8'h0, 8'h3b, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h2b, 8'h0, 8'h18, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h39, 8'h0, 8'h0, 8'h30, 8'h8c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h6c, 8'h0, 8'h0, 8'h38, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h96, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h70, 8'h26, 8'h0, 8'h2b, 8'h5d, 8'h83, 8'h8c, 8'h5d, 8'h1, 8'h0, 8'h44, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h55, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h0, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h69, 8'h96, 8'h98, 8'h9a, 8'h97, 8'h7d, 8'h34, 8'h0, 8'hf, 8'h65, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h3e, 8'h0, 8'h0, 8'h29, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h87, 8'h3d, 8'h12, 8'h2b, 8'h68, 8'h8d, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h7a, 8'h22, 8'h0, 8'h0, 8'h5c, 8'h95, 8'h9b, 8'h97, 8'h70, 8'h0, 8'h0, 8'h0, 8'h60, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8c, 8'h72, 8'h5f, 8'h60, 8'h65, 8'h6c, 8'h72, 8'h76, 8'h84, 8'h92, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h91, 8'h83, 8'h73, 8'h6f, 8'h6b, 8'h5c, 8'h21, 8'h0, 8'h0, 8'h49, 8'h5d, 8'hf, 8'h0, 8'h22, 8'h69, 8'h6d, 8'h48, 8'h4f, 8'h84, 8'h99, 8'h9a, 8'h9b, 8'h94, 8'h75, 8'h46, 8'h51, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h61, 8'h1a, 8'h0, 8'h0, 8'h14, 8'h4d, 8'h8f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8c, 8'h49, 8'h0, 8'h9, 8'h5e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6e, 8'h38, 8'h18, 8'h33, 8'h57, 8'h5e, 8'h42, 8'h14, 8'h0, 8'h15, 8'h45, 8'h74, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'hc, 8'h0, 8'h28, 8'h78, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h39, 8'h1e, 8'h20, 8'h42, 8'h7d, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3a, 8'h4, 8'h24, 8'h71, 8'h8c, 8'h97, 8'h99, 8'h8a, 8'h48, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h38, 8'h0, 8'h0, 8'h4d, 8'h94, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h71, 8'h0, 8'h0, 8'h2e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h73, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h20, 8'h6b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h68, 8'h0, 8'h0, 8'h2a, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h76, 8'h3, 8'h0, 8'h0, 8'h50, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7b, 8'h6e, 8'h7d, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h50, 8'h0, 8'h0, 8'h20, 8'h72, 8'h9b, 8'h9b, 8'h89, 8'h3b, 8'h0, 8'h0, 8'h16, 8'h80, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h8a, 8'h76, 8'h70, 8'h69, 8'h62, 8'h62, 8'h67, 8'h77, 8'h8b, 8'h96, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h96, 8'h95, 8'h88, 8'h70, 8'h46, 8'ha, 8'h0, 8'h2, 8'h4, 8'h0, 8'h0, 8'h57, 8'h8b, 8'h97, 8'h92, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h81, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h6d, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h33, 8'h42, 8'h46, 8'h58, 8'h7d, 8'h96, 8'h9b, 8'h9b, 8'h96, 8'h74, 8'hd, 8'h0, 8'h3c, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h50, 8'h0, 8'h0, 8'h0, 8'h4, 8'h9, 8'h0, 8'h0, 8'h23, 8'h5b, 8'h84, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6f, 8'h20, 8'h0, 8'h17, 8'h67, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h56, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h85, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h50, 8'ha, 8'he, 8'h6a, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h75, 8'h7, 8'h0, 8'h26, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h72, 8'h21, 8'h0, 8'h0, 8'h47, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h67, 8'h0, 8'h0, 8'h37, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h70, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h25, 8'h74, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'h28, 8'h0, 8'h0, 8'h4d, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h46, 8'h0, 8'h0, 8'h7, 8'h80, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7b, 8'h2f, 8'h0, 8'h0, 8'h43, 8'h94, 8'h9a, 8'h99, 8'h7a, 8'h1e, 8'h0, 8'h0, 8'h50, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h8c, 8'h83, 8'h7d, 8'h6d, 8'h5a, 8'h55, 8'h5f, 8'h77, 8'h90, 8'h93, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h96, 8'h92, 8'h8c, 8'h86, 8'h81, 8'h7f, 8'h7e, 8'h7e, 8'h7f, 8'h83, 8'h8a, 8'h91, 8'h97, 8'h98, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h91, 8'h70, 8'h4, 8'h0, 8'h0, 8'h0, 8'h13, 8'h69, 8'h83, 8'h8d, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h85, 8'h50, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h5f, 8'h90, 8'h9b, 8'h98, 8'h87, 8'h47, 8'h0, 8'h1c, 8'h6c, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h7b, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h42, 8'h7f, 8'h94, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h73, 8'h27, 8'h0, 8'h0, 8'h63, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6e, 8'h23, 8'h0, 8'h3b, 8'h2d, 8'h0, 8'h0, 8'h52, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h5f, 8'h9, 8'h0, 8'h41, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7e, 8'h18, 8'h0, 8'h32, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8a, 8'h4d, 8'h0, 8'h0, 8'h49, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h94, 8'h6c, 8'h12, 8'h0, 8'h0, 8'h0, 8'h51, 8'h87, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h70, 8'h0, 8'h0, 8'h8, 8'h83, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h7b, 8'hc, 8'h0, 8'h0, 8'h43, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h5f, 8'h0, 8'h0, 8'h1e, 8'h7c, 8'h9b, 8'h9b, 8'h91, 8'h55, 8'h0, 8'h0, 8'h0, 8'h5e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h95, 8'h84, 8'h5f, 8'h45, 8'h45, 8'h5f, 8'h84, 8'h91, 8'h93, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h88, 8'h80, 8'h7c, 8'h79, 8'h72, 8'h66, 8'h5a, 8'h4f, 8'h45, 8'h40, 8'h3e, 8'h3e, 8'h42, 8'h49, 8'h56, 8'h66, 8'h71, 8'h7b, 8'h86, 8'h8f, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h72, 8'h33, 8'h33, 8'h59, 8'h4e, 8'h44, 8'h4a, 8'h64, 8'h87, 8'h95, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h92, 8'h85, 8'h6c, 8'h40, 8'h39, 8'h3d, 8'h51, 8'h75, 8'h95, 8'h9b, 8'h91, 8'h5e, 8'h0, 8'h0, 8'h51, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h44, 8'h1b, 8'h76, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h82, 8'h33, 8'h0, 8'h4a, 8'h79, 8'h86, 8'h88, 8'h91, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h80, 8'h25, 8'h0, 8'h0, 8'h68, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h41, 8'h0, 8'h3e, 8'h7c, 8'h84, 8'h3a, 8'h0, 8'h0, 8'h5c, 8'h92, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h6a, 8'h0, 8'h0, 8'h3a, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h6a, 8'hb, 8'h25, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7d, 8'h30, 8'h0, 8'h7, 8'h62, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h6, 8'h58, 8'h8c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h46, 8'h0, 8'h0, 8'h10, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h57, 8'h0, 8'h0, 8'h0, 8'h64, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h3c, 8'h0, 8'h0, 8'h35, 8'h9a, 8'h9b, 8'h98, 8'h82, 8'h35, 8'h0, 8'h0, 8'h20, 8'h73, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7e, 8'h5d, 8'h4d, 8'h59, 8'h6f, 8'h7e, 8'h81, 8'h89, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h91, 8'h87, 8'h72, 8'h50, 8'h2d, 8'hf, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h25, 8'h52, 8'h7b, 8'h90, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h92, 8'h84, 8'h83, 8'h8e, 8'h88, 8'h82, 8'h7d, 8'h6b, 8'h51, 8'h4c, 8'h5d, 8'h82, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h86, 8'h84, 8'h85, 8'h8a, 8'h91, 8'h9a, 8'h98, 8'h82, 8'h35, 8'h0, 8'h10, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h44, 8'h0, 8'hf, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h41, 8'h0, 8'h36, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h2d, 8'h0, 8'h4, 8'h5e, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h58, 8'h10, 8'h5, 8'h76, 8'h95, 8'h98, 8'h7d, 8'h35, 8'h0, 8'h0, 8'h1d, 8'h58, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h85, 8'h43, 8'h0, 8'h35, 8'h7b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h71, 8'h8, 8'h0, 8'h47, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6b, 8'h18, 8'h0, 8'h2a, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h78, 8'h23, 8'h0, 8'h12, 8'h69, 8'h9b, 8'h94, 8'h6f, 8'h2e, 8'h0, 8'h0, 8'h0, 8'h13, 8'h5c, 8'h8a, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h76, 8'h1e, 8'h0, 8'h0, 8'h45, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h80, 8'h2f, 8'h0, 8'h0, 8'h15, 8'h6b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h94, 8'h9b, 8'h94, 8'h6d, 8'h14, 8'h0, 8'h0, 8'h2d, 8'h77, 8'h87, 8'h69, 8'h61, 8'h62, 8'h66, 8'h70, 8'h78, 8'h8a, 8'h97, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h94, 8'h85, 8'h68, 8'h45, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h53, 8'h79, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h99, 8'h96, 8'h86, 8'h75, 8'h6e, 8'h6b, 8'h65, 8'h61, 8'h69, 8'h80, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h8e, 8'h4b, 8'h0, 8'h0, 8'h50, 8'h88, 8'h9a, 8'h9b, 8'h96, 8'h6d, 8'h17, 8'h3, 8'h4b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h4c, 8'h0, 8'he, 8'h6c, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h62, 8'h0, 8'h2, 8'h48, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h32, 8'he, 8'h53, 8'h90, 8'h9b, 8'h99, 8'h95, 8'h7a, 8'h2c, 8'h0, 8'h0, 8'h27, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h53, 8'h0, 8'h0, 8'h62, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h66, 8'h13, 8'h0, 8'h37, 8'h78, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h3c, 8'hf, 8'h27, 8'h73, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h77, 8'h24, 8'h0, 8'h14, 8'h68, 8'h83, 8'h52, 8'h18, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h67, 8'h8d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h57, 8'h0, 8'h0, 8'h0, 8'h63, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h60, 8'ha, 8'h0, 8'h0, 8'h35, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h2e, 8'h0, 8'h0, 8'h26, 8'h88, 8'h99, 8'h9b, 8'h90, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h33, 8'h6b, 8'h62, 8'h61, 8'h6f, 8'h86, 8'h95, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h80, 8'h66, 8'h43, 8'he, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h6d, 8'h8e, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h94, 8'h89, 8'h72, 8'h5e, 8'h5e, 8'h65, 8'h6f, 8'h78, 8'h89, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h7a, 8'h1d, 8'h0, 8'hb, 8'h7c, 8'h99, 8'h9b, 8'h9a, 8'h88, 8'h32, 8'h0, 8'h27, 8'h82, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h5d, 8'h0, 8'h0, 8'h5f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h6a, 8'h1a, 8'h0, 8'h32, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h52, 8'h13, 8'h27, 8'h8b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h86, 8'h37, 8'h0, 8'h0, 8'h45, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h35, 8'h0, 8'h0, 8'h6f, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h65, 8'h1c, 8'h0, 8'h33, 8'h77, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h40, 8'h13, 8'h25, 8'h6a, 8'h94, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h33, 8'h0, 8'ha, 8'h47, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h82, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h40, 8'h0, 8'h0, 8'h38, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h50, 8'h0, 8'h0, 8'h0, 8'h51, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h76, 8'h16, 8'h0, 8'h0, 8'h6e, 8'h94, 8'h99, 8'h90, 8'h6e, 8'h1b, 8'h0, 8'h0, 8'h14, 8'h63, 8'h88, 8'h93, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8c, 8'h71, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h6a, 8'h90, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h92, 8'h85, 8'h64, 8'h53, 8'h56, 8'h6c, 8'h86, 8'h88, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h4c, 8'h0, 8'h0, 8'h54, 8'h8e, 8'h9b, 8'h9a, 8'h92, 8'h62, 8'h0, 8'h7, 8'h57, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6e, 8'h17, 8'h0, 8'h5b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h72, 8'h27, 8'h0, 8'he, 8'h64, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h64, 8'h10, 8'hc, 8'h50, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h8b, 8'h57, 8'h0, 8'h0, 8'h48, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h41, 8'h0, 8'h0, 8'h57, 8'h8c, 8'h9b, 8'h9b, 8'h94, 8'h6a, 8'h1b, 8'h0, 8'h22, 8'h7f, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h57, 8'h0, 8'h1b, 8'h64, 8'h96, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h59, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6e, 8'h11, 8'h0, 8'h0, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h3a, 8'h0, 8'h0, 8'h16, 8'h83, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h55, 8'h0, 8'h0, 8'h40, 8'h80, 8'h90, 8'h73, 8'h43, 8'h35, 8'h39, 8'h57, 8'h7f, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h92, 8'h86, 8'h68, 8'h3a, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h62, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h8f, 8'h82, 8'h65, 8'h43, 8'h4a, 8'h73, 8'h8f, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h79, 8'h0, 8'h0, 8'h11, 8'h93, 8'h9a, 8'h9a, 8'h96, 8'h70, 8'h17, 8'h0, 8'h49, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h69, 8'h11, 8'h0, 8'h5b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h83, 8'h2c, 8'h0, 8'h0, 8'h69, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6a, 8'h0, 8'h0, 8'h47, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h54, 8'h0, 8'h0, 8'h51, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h80, 8'h3d, 8'h0, 8'h0, 8'h58, 8'h96, 8'h96, 8'h79, 8'he, 8'h0, 8'h1f, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h62, 8'h0, 8'h0, 8'h52, 8'h95, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h57, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h6c, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h56, 8'h0, 8'h0, 8'h2d, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h70, 8'h2, 8'h0, 8'h0, 8'h25, 8'h8d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h4f, 8'h1b, 8'h4f, 8'h53, 8'h54, 8'h63, 8'h78, 8'h7c, 8'h81, 8'h8c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h98, 8'h9b, 8'h99, 8'h9a, 8'h96, 8'h8c, 8'h73, 8'h54, 8'h36, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h6b, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8b, 8'h7c, 8'h78, 8'h60, 8'h52, 8'h5a, 8'h77, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h81, 8'h27, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h52, 8'h0, 8'h13, 8'h6a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h53, 8'h0, 8'h0, 8'h64, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h37, 8'h0, 8'h0, 8'h65, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h5c, 8'h5, 8'h0, 8'h47, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h51, 8'h4, 8'h0, 8'h4e, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7d, 8'h3a, 8'h0, 8'h0, 8'h7, 8'h12, 8'h0, 8'h0, 8'h24, 8'h77, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h93, 8'h65, 8'h15, 8'h0, 8'h49, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h47, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h47, 8'h7c, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h78, 8'h5, 8'h0, 8'h0, 8'h56, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h49, 8'h0, 8'h0, 8'h0, 8'h45, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h80, 8'h54, 8'h36, 8'h58, 8'h67, 8'h70, 8'h7f, 8'h94, 8'h98, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h77, 8'h92, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h8f, 8'h6d, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h7d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h92, 8'h7c, 8'h6c, 8'h65, 8'h61, 8'h64, 8'h6d, 8'h85, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h56, 8'h0, 8'h0, 8'h34, 8'h87, 8'h9a, 8'h9a, 8'h94, 8'h69, 8'h17, 8'h0, 8'h4d, 8'h87, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8a, 8'h3e, 8'h0, 8'h32, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h55, 8'h1, 8'h0, 8'h45, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h7d, 8'h30, 8'h0, 8'h3f, 8'h81, 8'h98, 8'h9b, 8'h9b, 8'h8d, 8'h53, 8'hf, 8'h1, 8'h42, 8'h86, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7f, 8'h43, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h24, 8'h6d, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h61, 8'h1d, 8'h0, 8'h31, 8'h7b, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h5f, 8'h17, 8'h18, 8'h44, 8'h79, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h45, 8'h0, 8'h0, 8'h15, 8'h84, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h81, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h58, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h7f, 8'h75, 8'h69, 8'h5b, 8'h5a, 8'h70, 8'h8b, 8'h96, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h91, 8'h6e, 8'h27, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'ha, 8'h63, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h95, 8'h88, 8'h6f, 8'h5f, 8'h5f, 8'h6a, 8'h78, 8'h7e, 8'h93, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h6b, 8'h12, 8'h0, 8'h18, 8'h6c, 8'h99, 8'h9b, 8'h98, 8'h7f, 8'h36, 8'h0, 8'h17, 8'h7c, 8'h99, 8'h9a, 8'h9b, 8'h92, 8'h6f, 8'h5e, 8'h74, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h5f, 8'h13, 8'h0, 8'h63, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h75, 8'h16, 8'h0, 8'h2b, 8'h80, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h76, 8'h20, 8'h0, 8'h4e, 8'h82, 8'h98, 8'h99, 8'h8e, 8'h5c, 8'h11, 8'h6, 8'h3d, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8d, 8'h6f, 8'h34, 8'h0, 8'h1c, 8'h6c, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h6a, 8'h21, 8'h0, 8'h22, 8'h78, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h88, 8'h8a, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7b, 8'he, 8'h0, 8'h0, 8'h4d, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h73, 8'h23, 8'h0, 8'h0, 8'h15, 8'h68, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8f, 8'h88, 8'h7a, 8'h57, 8'h51, 8'h66, 8'h83, 8'h93, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h9b, 8'h99, 8'h8b, 8'h66, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h7d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h97, 8'h91, 8'h82, 8'h65, 8'h4f, 8'h5a, 8'h79, 8'h88, 8'h91, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h3b, 8'h0, 8'h0, 8'h56, 8'h96, 8'h9b, 8'h9b, 8'h8f, 8'h57, 8'hc, 8'h3, 8'h6a, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h8a, 8'h3c, 8'h4, 8'h20, 8'h79, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8f, 8'h78, 8'h57, 8'h17, 8'h0, 8'h1d, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h3d, 8'h0, 8'h14, 8'h65, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h82, 8'h38, 8'h0, 8'h3, 8'h4a, 8'h71, 8'h7d, 8'h62, 8'hf, 8'h0, 8'h3c, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h90, 8'h86, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h81, 8'h6e, 8'h83, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h29, 8'h0, 8'h1c, 8'h6e, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h67, 8'h12, 8'h0, 8'h0, 8'h38, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8a, 8'h5e, 8'h41, 8'h50, 8'h7d, 8'h8d, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h8a, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h5c, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h93, 8'h8d, 8'h7d, 8'h50, 8'h47, 8'h63, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h65, 8'hd, 8'h0, 8'h1e, 8'h76, 8'h9b, 8'h9b, 8'h9a, 8'h7e, 8'h13, 8'h0, 8'h33, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h71, 8'h0, 8'h0, 8'h4, 8'h7a, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h56, 8'h0, 8'h0, 8'h0, 8'h23, 8'h88, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h4e, 8'h0, 8'h0, 8'h52, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h4, 8'h1, 8'h0, 8'h3c, 8'h81, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h5f, 8'h2c, 8'h69, 8'h99, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h54, 8'h0, 8'h1b, 8'h66, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'h33, 8'h0, 8'h0, 8'hd, 8'h6a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8c, 8'h51, 8'h0, 8'h0, 8'h0, 8'h49, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h7c, 8'h58, 8'h58, 8'h6a, 8'h7a, 8'h81, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h99, 8'h8d, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h86, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h80, 8'h76, 8'h68, 8'h55, 8'h59, 8'h7b, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h28, 8'h0, 8'h0, 8'h62, 8'h91, 8'h9b, 8'h99, 8'h82, 8'h26, 8'h0, 8'h1f, 8'h7e, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h30, 8'h0, 8'h0, 8'h0, 8'h16, 8'h44, 8'h67, 8'h74, 8'h70, 8'h3b, 8'h13, 8'h0, 8'h0, 8'h0, 8'h25, 8'h53, 8'h78, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h4f, 8'h0, 8'h0, 8'h45, 8'h84, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h86, 8'h62, 8'h44, 8'h2, 8'h0, 8'h0, 8'h2d, 8'h75, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h4a, 8'h3, 8'h27, 8'h40, 8'h2d, 8'h1f, 8'h65, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h58, 8'h0, 8'h0, 8'h4b, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h6b, 8'h17, 8'h0, 8'h0, 8'h34, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h31, 8'h0, 8'h0, 8'h6, 8'h68, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h73, 8'h64, 8'h64, 8'h6a, 8'h71, 8'h87, 8'h96, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h31, 8'h42, 8'h46, 8'h40, 8'h32, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h7d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h95, 8'h83, 8'h6e, 8'h67, 8'h63, 8'h66, 8'h75, 8'h8a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h45, 8'h0, 8'h0, 8'h26, 8'h87, 8'h99, 8'h9a, 8'h93, 8'h65, 8'h0, 8'h12, 8'h5f, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h6c, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9, 8'h7, 8'h0, 8'h0, 8'h0, 8'h20, 8'h44, 8'h74, 8'h8f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h5d, 8'hf, 8'h0, 8'h30, 8'h7e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h86, 8'h58, 8'h30, 8'h3f, 8'h73, 8'h91, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h84, 8'h4a, 8'h9, 8'hd, 8'h59, 8'h5f, 8'h26, 8'h0, 8'hd, 8'h51, 8'h85, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h59, 8'h5, 8'h0, 8'h35, 8'h79, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h5b, 8'h0, 8'h0, 8'h0, 8'h53, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h74, 8'h10, 8'h0, 8'h0, 8'h24, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h88, 8'h77, 8'h6c, 8'h5f, 8'h5e, 8'h70, 8'h92, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h64, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h3a, 8'h4c, 8'h5f, 8'h6f, 8'h7e, 8'h8b, 8'h90, 8'h91, 8'h8e, 8'h84, 8'h70, 8'h53, 8'h15, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h70, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h96, 8'h8c, 8'h6e, 8'h5e, 8'h60, 8'h6c, 8'h7a, 8'h88, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6e, 8'h8, 8'h0, 8'he, 8'h70, 8'h94, 8'h9b, 8'h97, 8'h7b, 8'h32, 8'h0, 8'h44, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h79, 8'h41, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h16, 8'h41, 8'h78, 8'h8e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h78, 8'h21, 8'h0, 8'h1b, 8'h7f, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h85, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h8e, 8'h91, 8'h97, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h4f, 8'h13, 8'h8, 8'h51, 8'h87, 8'h8c, 8'h5d, 8'h16, 8'h0, 8'hf, 8'h60, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5e, 8'he, 8'h0, 8'h18, 8'h77, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h4d, 8'h0, 8'h0, 8'h1d, 8'h86, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h93, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h69, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8d, 8'h7e, 8'h65, 8'h4c, 8'h59, 8'h7c, 8'h93, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7c, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h30, 8'h60, 8'h7e, 8'h89, 8'h91, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h96, 8'h92, 8'h7e, 8'h69, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h5a, 8'h8a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h94, 8'h92, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h8f, 8'h8e, 8'h8f, 8'h8f, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h8e, 8'h79, 8'h59, 8'h4e, 8'h65, 8'h7f, 8'h8e, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h84, 8'h37, 8'h0, 8'h0, 8'h50, 8'h97, 8'h9b, 8'h99, 8'h8c, 8'h51, 8'h0, 8'h0, 8'h61, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h85, 8'h77, 8'h5a, 8'h48, 8'h4e, 8'h62, 8'h7c, 8'h8a, 8'h91, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h46, 8'h0, 8'h7, 8'h5c, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h65, 8'h49, 8'h5a, 8'h89, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8d, 8'h54, 8'ha, 8'h6, 8'h4a, 8'h92, 8'h99, 8'h9a, 8'h91, 8'h6d, 8'h1f, 8'h0, 8'h2d, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h6c, 8'hd, 8'h0, 8'h14, 8'h7f, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h76, 8'h0, 8'h0, 8'h0, 8'h44, 8'h94, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h82, 8'h25, 8'h0, 8'h0, 8'h13, 8'h74, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h7a, 8'h56, 8'h48, 8'h61, 8'h89, 8'h8f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h82, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h56, 8'h77, 8'h8d, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h87, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h80, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h93, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h77, 8'h54, 8'h36, 8'h31, 8'h37, 8'h3a, 8'h51, 8'h7c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8f, 8'h83, 8'h5f, 8'h4d, 8'h58, 8'h7e, 8'h98, 8'h9b, 8'h9b, 8'h97, 8'h65, 8'h0, 8'h0, 8'h35, 8'h90, 8'h9b, 8'h9a, 8'h95, 8'h72, 8'h21, 8'h0, 8'h4a, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h92, 8'h8f, 8'h91, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h62, 8'h0, 8'h0, 8'h3e, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h97, 8'h74, 8'h0, 8'h0, 8'h0, 8'h30, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h90, 8'h60, 8'h0, 8'h1, 8'h49, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h67, 8'h0, 8'h0, 8'h3e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h78, 8'h5, 8'h0, 8'h1a, 8'h77, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h49, 8'h0, 8'h0, 8'hc, 8'h8b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h65, 8'hb, 8'h0, 8'h0, 8'h3d, 8'h82, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h78, 8'h58, 8'h5b, 8'h6c, 8'h7b, 8'h87, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h53, 8'h72, 8'h88, 8'h95, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h76, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h7f, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h76, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h87, 8'h78, 8'h69, 8'h5a, 8'h5a, 8'h76, 8'h8c, 8'h82, 8'h3c, 8'h0, 8'h1a, 8'h6e, 8'h9a, 8'h9b, 8'h9b, 8'h8b, 8'h40, 8'h0, 8'h2, 8'h74, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h63, 8'h4, 8'h0, 8'h34, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h6b, 8'h9, 8'h0, 8'h11, 8'hd, 8'h0, 8'h2b, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h53, 8'h0, 8'h0, 8'h42, 8'h85, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h64, 8'h0, 8'ha, 8'h5f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h61, 8'h1, 8'h0, 8'h1b, 8'h65, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h76, 8'hc, 8'h0, 8'h0, 8'h50, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h89, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h53, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h77, 8'h68, 8'h65, 8'h67, 8'h73, 8'h8b, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7a, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h64, 8'h8b, 8'h95, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h48, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h16, 8'h6e, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h64, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h83, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h94, 8'h89, 8'h70, 8'h65, 8'h63, 8'h5f, 8'h40, 8'h0, 8'h0, 8'h4c, 8'h8e, 8'h9b, 8'h9b, 8'h96, 8'h70, 8'h1b, 8'h0, 8'h4b, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6a, 8'h1c, 8'h0, 8'h1b, 8'h6f, 8'h99, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h72, 8'h2f, 8'h0, 8'h1d, 8'h5c, 8'h56, 8'hc, 8'h0, 8'h33, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8b, 8'h53, 8'h6, 8'h0, 8'h3b, 8'h7c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h73, 8'h1d, 8'h0, 8'h3b, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5c, 8'hb, 8'h0, 8'he, 8'h5d, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h3d, 8'h0, 8'h0, 8'h5, 8'h6f, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7e, 8'h38, 8'h0, 8'h0, 8'h13, 8'h6d, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8f, 8'h7a, 8'h72, 8'h5f, 8'h5f, 8'h72, 8'h94, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h50, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h74, 8'h96, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h66, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h6b, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h5e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h52, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h96, 8'h8d, 8'h70, 8'h52, 8'h15, 8'h0, 8'h0, 8'h5f, 8'h96, 8'h9b, 8'h9b, 8'h8a, 8'h42, 8'h3, 8'h19, 8'h89, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h71, 8'h2a, 8'h0, 8'h0, 8'h62, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h60, 8'h2c, 8'h0, 8'h0, 8'h5f, 8'h8e, 8'h8d, 8'h5b, 8'h0, 8'h0, 8'h50, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h68, 8'h14, 8'h0, 8'h2c, 8'h7f, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h78, 8'h2f, 8'h0, 8'h1b, 8'h69, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h65, 8'h12, 8'h0, 8'h0, 8'h5a, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7a, 8'h1f, 8'h0, 8'h0, 8'h44, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h72, 8'hd, 8'h0, 8'h0, 8'h22, 8'h90, 8'h98, 8'h93, 8'h8a, 8'h71, 8'h4a, 8'h57, 8'h7e, 8'h92, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h74, 8'h15, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h79, 8'h97, 8'h9a, 8'h9a, 8'h99, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h6a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'he, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h84, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h83, 8'h35, 8'h0, 8'h4, 8'h5c, 8'h89, 8'h94, 8'h93, 8'h6a, 8'h6, 8'h0, 8'h48, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h33, 8'h0, 8'h0, 8'h52, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h1b, 8'h0, 8'h0, 8'h3a, 8'h84, 8'h9a, 8'h9a, 8'h88, 8'h49, 8'h0, 8'h38, 8'h8d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h3e, 8'h0, 8'h0, 8'h77, 8'h8d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h3b, 8'h0, 8'h0, 8'h6a, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h77, 8'h13, 8'h0, 8'h0, 8'h57, 8'h8a, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h53, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h61, 8'h0, 8'h0, 8'h0, 8'h49, 8'h82, 8'h64, 8'h4d, 8'h5e, 8'h84, 8'h8b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h7f, 8'h97, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h6e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h6b, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h32, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h80, 8'h64, 8'h70, 8'h54, 8'h4d, 8'h66, 8'h74, 8'hf, 8'h0, 8'h30, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h6e, 8'h3, 8'h0, 8'h45, 8'h8e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6a, 8'hf, 8'h22, 8'h7a, 8'h88, 8'h97, 8'h9b, 8'h97, 8'h7c, 8'h2a, 8'h0, 8'h3a, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h63, 8'h5, 8'h0, 8'h0, 8'h4b, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h65, 8'h12, 8'h0, 8'h66, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h37, 8'h0, 8'h0, 8'h49, 8'h8e, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7e, 8'h33, 8'h0, 8'h0, 8'h2a, 8'h7e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h36, 8'h0, 8'h0, 8'h0, 8'h46, 8'h65, 8'h73, 8'h84, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h77, 8'h16, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h40, 8'h85, 8'h98, 8'h97, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h69, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h6c, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h92, 8'h93, 8'h7e, 8'h73, 8'h64, 8'h36, 8'h0, 8'h13, 8'h64, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h71, 8'ha, 8'h0, 8'h24, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h74, 8'h1b, 8'hb, 8'h4c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h60, 8'h0, 8'h14, 8'h62, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h5b, 8'h1b, 8'h0, 8'h0, 8'h14, 8'h4f, 8'h87, 8'h9a, 8'h85, 8'h2c, 8'h0, 8'h23, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h5d, 8'h0, 8'h0, 8'h2b, 8'h82, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h68, 8'h0, 8'h0, 8'h0, 8'h21, 8'h59, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h5e, 8'h4, 8'h0, 8'h0, 8'h21, 8'h6f, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h89, 8'h99, 8'h96, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h56, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h74, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h2e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h98, 8'h8f, 8'h60, 8'h4, 8'h0, 8'h20, 8'h62, 8'h86, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h96, 8'h6e, 8'h1c, 8'h0, 8'h8, 8'h5d, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h77, 8'h2a, 8'h0, 8'h30, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6d, 8'h21, 8'h0, 8'h4b, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8e, 8'h6e, 8'h37, 8'h12, 8'h0, 8'h0, 8'h36, 8'h5f, 8'h3e, 8'h0, 8'ha, 8'h64, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h61, 8'h9, 8'h0, 8'h19, 8'h69, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8d, 8'h54, 8'h0, 8'h0, 8'h0, 8'h9, 8'h89, 8'h9a, 8'h9b, 8'h97, 8'h8f, 8'h7b, 8'h5f, 8'h2b, 8'h0, 8'h0, 8'h33, 8'h7d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7f, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5e, 8'h8f, 8'h9a, 8'h98, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h36, 8'h7c, 8'h97, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h74, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h60, 8'hc, 8'h6, 8'h38, 8'h56, 8'h6a, 8'h81, 8'h8f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h82, 8'h37, 8'h0, 8'h0, 8'h56, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h3e, 8'h0, 8'h20, 8'h6d, 8'h97, 8'h9b, 8'h9b, 8'h98, 8'h7b, 8'h34, 8'h0, 8'h1e, 8'h78, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h8b, 8'h6a, 8'h27, 8'h0, 8'h0, 8'h4, 8'h0, 8'h0, 8'h43, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h66, 8'h15, 8'h0, 8'h1, 8'h62, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h71, 8'h92, 8'h94, 8'h89, 8'h6c, 8'h4a, 8'h59, 8'h72, 8'h6c, 8'h4e, 8'h7a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h68, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h71, 8'h93, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h1e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4f, 8'h86, 8'h99, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7f, 8'h60, 8'h79, 8'h87, 8'h78, 8'h57, 8'h4c, 8'h6f, 8'h89, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h5a, 8'hb, 8'h0, 8'h61, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h4f, 8'h5, 8'h0, 8'h6d, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h48, 8'h4, 8'h8, 8'h7a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h85, 8'h84, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h87, 8'h5b, 8'h17, 8'h0, 8'h0, 8'h36, 8'h83, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'h11, 8'h0, 8'h0, 8'h63, 8'h8f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h7e, 8'h3c, 8'h0, 8'h0, 8'h4, 8'h66, 8'h6a, 8'h4f, 8'h59, 8'h80, 8'h8b, 8'h93, 8'h95, 8'h8c, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h5a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h7c, 8'h97, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h67, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h65, 8'h8f, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h79, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h90, 8'h98, 8'h99, 8'h94, 8'h8b, 8'h7a, 8'h59, 8'h51, 8'h71, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h67, 8'h14, 8'h0, 8'h15, 8'h82, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h48, 8'h7, 8'hd, 8'h6b, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h8c, 8'h46, 8'h4, 8'hd, 8'h5e, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h7f, 8'h20, 8'h0, 8'h35, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h67, 8'h26, 8'h15, 8'h60, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h7c, 8'hc, 8'h0, 8'h0, 8'h63, 8'h8e, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h7d, 8'h5a, 8'h20, 8'h0, 8'h10, 8'h4d, 8'h71, 8'h7e, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h94, 8'h49, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h82, 8'h98, 8'h9b, 8'h99, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h74, 8'h95, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h7d, 8'h71, 8'h65, 8'h60, 8'h70, 8'h92, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h6d, 8'h18, 8'h0, 8'h14, 8'h68, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h2a, 8'h0, 8'h0, 8'h5a, 8'h86, 8'h97, 8'h99, 8'h8a, 8'h54, 8'ha, 8'h14, 8'h51, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8f, 8'h69, 8'h20, 8'h0, 8'h0, 8'h0, 8'h40, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h77, 8'h6a, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h7c, 8'h22, 8'h0, 8'h0, 8'h54, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h75, 8'h45, 8'h0, 8'h0, 8'h4b, 8'h90, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h90, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h63, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h85, 8'h99, 8'h9b, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h29, 8'h7c, 8'h97, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h69, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h91, 8'h7b, 8'h63, 8'h63, 8'h6f, 8'h7c, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h67, 8'h1d, 8'h0, 8'h11, 8'h5e, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h4f, 8'hd, 8'h0, 8'h12, 8'h31, 8'h4c, 8'h63, 8'h57, 8'hf, 8'hd, 8'h4a, 8'h83, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h68, 8'h1b, 8'h0, 8'h27, 8'h1b, 8'h0, 8'h0, 8'h7a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h84, 8'h46, 8'h0, 8'h0, 8'h3d, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h88, 8'h84, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h85, 8'h73, 8'h5e, 8'h50, 8'h4d, 8'h36, 8'h67, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h98, 8'h88, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h77, 8'h69, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h38, 8'h89, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h83, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h8e, 8'h7b, 8'h59, 8'h5d, 8'h72, 8'h89, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6c, 8'h1d, 8'h0, 8'h7, 8'h5a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h5a, 8'h22, 8'h6, 8'h0, 8'h0, 8'he, 8'h16, 8'h0, 8'h45, 8'h7f, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h76, 8'h27, 8'h0, 8'h2f, 8'h72, 8'h6b, 8'h1c, 8'h0, 8'h52, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h57, 8'h2, 8'h0, 8'h20, 8'h6f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h4e, 8'h41, 8'h65, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h97, 8'h86, 8'h54, 8'h4b, 8'h6b, 8'h92, 8'h91, 8'h90, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h91, 8'h61, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h79, 8'h8d, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h83, 8'h29, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4b, 8'h89, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8b, 8'h6a, 8'h4f, 8'h59, 8'h88, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h85, 8'h31, 8'h0, 8'h0, 8'h5f, 8'h93, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8c, 8'h85, 8'h66, 8'ha, 8'h0, 8'h0, 8'h38, 8'h80, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h84, 8'h2f, 8'h0, 8'h0, 8'h7b, 8'h96, 8'h8c, 8'h41, 8'h0, 8'h0, 8'h61, 8'h8e, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h65, 8'h12, 8'h0, 8'h0, 8'h65, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h82, 8'h5d, 8'h52, 8'h6f, 8'h80, 8'h8f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h87, 8'h37, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h73, 8'h96, 8'h8a, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h16, 8'h67, 8'h90, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8d, 8'h84, 8'h6e, 8'h4f, 8'h5d, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h3e, 8'h0, 8'h0, 8'h51, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h91, 8'h71, 8'h54, 8'h58, 8'h82, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h36, 8'h0, 8'h0, 8'h58, 8'h92, 8'h9b, 8'h95, 8'h70, 8'h1d, 8'h0, 8'h0, 8'h2, 8'h3a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h62, 8'hf, 8'h0, 8'h0, 8'h63, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h86, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h71, 8'h5e, 8'h62, 8'h73, 8'h8d, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9a, 8'h99, 8'h80, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h6e, 8'h96, 8'h9a, 8'h83, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h90, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h84, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h71, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h8b, 8'h6f, 8'h61, 8'h61, 8'h72, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h40, 8'h0, 8'h0, 8'h1b, 8'h82, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8f, 8'h6b, 8'h48, 8'h70, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h8c, 8'h8b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h44, 8'h0, 8'h0, 8'h40, 8'h89, 8'h9a, 8'h9b, 8'h98, 8'h8f, 8'h65, 8'h16, 8'h0, 8'h0, 8'h1c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h65, 8'hf, 8'h0, 8'h0, 8'h56, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h53, 8'h2b, 8'h49, 8'h77, 8'h92, 8'h99, 8'h92, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h77, 8'h6b, 8'h64, 8'h6b, 8'h80, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h7a, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h92, 8'h9b, 8'h99, 8'h7e, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h6f, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h90, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h72, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h80, 8'h68, 8'h62, 8'h69, 8'h7a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h60, 8'h0, 8'h0, 8'hf, 8'h5f, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h76, 8'h6a, 8'h42, 8'h0, 8'h22, 8'h5d, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h64, 8'h2, 8'h0, 8'h32, 8'h7a, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h4d, 8'h1, 8'h0, 8'h38, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h6d, 8'h17, 8'h0, 8'h0, 8'h4e, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h66, 8'hc, 8'h0, 8'h0, 8'h2d, 8'h67, 8'h8a, 8'h8e, 8'h54, 8'h0, 8'h0, 8'h4, 8'h0, 8'h0, 8'h2, 8'h55, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h8a, 8'h74, 8'h54, 8'h59, 8'h7d, 8'h95, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h80, 8'h39, 8'h0, 8'h0, 8'h0, 8'h37, 8'h88, 8'h9a, 8'h9b, 8'h99, 8'h7a, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h7a, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h6f, 8'h96, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h74, 8'h53, 8'h58, 8'h7b, 8'h8d, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h75, 8'h1c, 8'h0, 8'h7, 8'h58, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h67, 8'h2f, 8'h42, 8'h48, 8'h0, 8'h0, 8'h1c, 8'h63, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h78, 8'h2c, 8'h0, 8'h26, 8'h71, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h84, 8'h41, 8'h5, 8'h20, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h78, 8'h2d, 8'h0, 8'h0, 8'h4f, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h65, 8'h8, 8'h0, 8'h0, 8'h0, 8'h1, 8'h50, 8'h89, 8'h50, 8'h0, 8'h0, 8'h43, 8'h3b, 8'h0, 8'h0, 8'hf, 8'h6a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h82, 8'h5e, 8'h4c, 8'h70, 8'h8b, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h98, 8'h8d, 8'h7c, 8'h60, 8'h44, 8'h52, 8'h81, 8'h98, 8'h9b, 8'h9b, 8'h98, 8'h7b, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h84, 8'h40, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8c, 8'h75, 8'h4e, 8'h5c, 8'h7f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8b, 8'h4a, 8'h0, 8'h0, 8'h47, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6c, 8'h0, 8'h0, 8'h3b, 8'h8d, 8'h79, 8'h3e, 8'h2, 8'h32, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h86, 8'h37, 8'h0, 8'h0, 8'h65, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h58, 8'h0, 8'h1f, 8'h66, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h38, 8'h0, 8'h0, 8'h57, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h80, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h13, 8'h0, 8'h9, 8'h62, 8'h78, 8'h23, 8'h0, 8'h0, 8'h19, 8'h84, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h63, 8'h55, 8'h68, 8'h82, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9b, 8'h99, 8'h96, 8'h94, 8'h90, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h77, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h8d, 8'h9a, 8'h97, 8'h8d, 8'h8e, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8f, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h6d, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h7b, 8'h60, 8'h51, 8'h65, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h45, 8'h0, 8'h0, 8'h38, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h63, 8'h7, 8'h0, 8'h2c, 8'h75, 8'h9b, 8'h97, 8'h70, 8'h8, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h85, 8'h31, 8'h0, 8'h0, 8'h55, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h4c, 8'h1, 8'h1c, 8'h62, 8'h8f, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h39, 8'h0, 8'h0, 8'h3a, 8'h82, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h2b, 8'h0, 8'h0, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h78, 8'h92, 8'h64, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h91, 8'h99, 8'h8f, 8'h78, 8'h61, 8'h63, 8'h6f, 8'h85, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h76, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h8c, 8'h91, 8'h6d, 8'h35, 8'h2c, 8'h59, 8'h85, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h74, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h83, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h81, 8'h6e, 8'h65, 8'h66, 8'h79, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h45, 8'h0, 8'h0, 8'h27, 8'h75, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h69, 8'h1f, 8'h0, 8'h2a, 8'h70, 8'h94, 8'h9b, 8'h9b, 8'h80, 8'h17, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h83, 8'h47, 8'hf, 8'h13, 8'h60, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3a, 8'h0, 8'h0, 8'hd, 8'h77, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8c, 8'h3f, 8'h0, 8'h0, 8'h42, 8'h3c, 8'hd, 8'h0, 8'h0, 8'h0, 8'h47, 8'h8c, 8'h9a, 8'h88, 8'h3c, 8'h0, 8'h0, 8'h20, 8'h7a, 8'h7e, 8'h6d, 8'h61, 8'h62, 8'h7f, 8'h8f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h75, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h86, 8'h75, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h8d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h32, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h29, 8'h72, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h27, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h67, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h92, 8'h81, 8'h61, 8'h60, 8'h6f, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h6a, 8'h9, 8'h0, 8'h19, 8'h74, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h39, 8'h0, 8'hc, 8'h71, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h7f, 8'h1a, 8'hc, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h64, 8'h26, 8'h0, 8'h0, 8'h0, 8'h38, 8'h7b, 8'h99, 8'h99, 8'h87, 8'h48, 8'hc, 8'he, 8'h58, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h52, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h7d, 8'h67, 8'h70, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h5c, 8'h0, 8'h0, 8'h46, 8'h7f, 8'h7f, 8'h60, 8'h3f, 8'h5b, 8'h81, 8'h98, 8'h9b, 8'h99, 8'h7f, 8'h29, 8'h0, 8'h0, 8'h50, 8'h57, 8'h54, 8'h6c, 8'h93, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h74, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h72, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h6d, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h8b, 8'h6a, 8'h57, 8'h66, 8'h8a, 8'h93, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7d, 8'h2f, 8'h0, 8'h4, 8'h68, 8'h94, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h65, 8'h11, 8'h0, 8'h54, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h63, 8'h11, 8'h34, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h89, 8'h79, 8'h4e, 8'h0, 8'h0, 8'h34, 8'h80, 8'h8c, 8'h57, 8'h3, 8'h6, 8'h4d, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h7e, 8'h1b, 8'h0, 8'h0, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6a, 8'h14, 8'h0, 8'h3b, 8'h80, 8'h99, 8'h96, 8'h91, 8'h94, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h2f, 8'h0, 8'h17, 8'h59, 8'h83, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h73, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h29, 8'h38, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h76, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h79, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h91, 8'h83, 8'h74, 8'h6b, 8'h77, 8'h85, 8'h90, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'he, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h43, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h84, 8'h65, 8'h46, 8'h6e, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h84, 8'h40, 8'h0, 8'h0, 8'h2f, 8'h97, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h80, 8'h14, 8'h0, 8'h26, 8'h94, 8'h9b, 8'h99, 8'h9b, 8'h9a, 8'h76, 8'h7, 8'h2, 8'h4d, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8e, 8'h59, 8'h0, 8'h0, 8'h26, 8'h64, 8'h0, 8'h0, 8'h48, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h35, 8'h0, 8'h0, 8'h3e, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h74, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h7d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h92, 8'h60, 8'h3, 8'h0, 8'h34, 8'h7f, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h72, 8'h3f, 8'h29, 8'h67, 8'h87, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h71, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h83, 8'h99, 8'h9b, 8'h9b, 8'h99, 8'h73, 8'hc, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h5e, 8'h8d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h81, 8'h5e, 8'h36, 8'h7, 8'h0, 8'h0, 8'h20, 8'h4b, 8'h79, 8'h93, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h76, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h6f, 8'h56, 8'h5e, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h80, 8'h40, 8'h0, 8'h0, 8'h2a, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h40, 8'h0, 8'h1a, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h68, 8'hd, 8'h0, 8'h42, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h7c, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h3e, 8'h0, 8'h0, 8'h31, 8'h7c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h77, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h56, 8'h28, 8'h29, 8'h26, 8'h25, 8'h8, 8'h0, 8'h0, 8'h4f, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h70, 8'h5e, 8'h60, 8'h73, 8'h92, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5f, 8'h93, 8'h9a, 8'h9a, 8'h8a, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h49, 8'h82, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h64, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h71, 8'h8f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h72, 8'h66, 8'h64, 8'h75, 8'h90, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h4c, 8'h0, 8'h0, 8'h26, 8'h72, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6f, 8'h0, 8'h0, 8'h1c, 8'h76, 8'h9b, 8'h9a, 8'h92, 8'h65, 8'h1d, 8'h0, 8'h3d, 8'h7c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'h4e, 8'h3f, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h87, 8'h4c, 8'h3, 8'h0, 8'h0, 8'h57, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8b, 8'h42, 8'h0, 8'h0, 8'hc, 8'h70, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h75, 8'h2d, 8'h0, 8'h8, 8'h4d, 8'h55, 8'h5, 8'hc, 8'h51, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h9a, 8'h99, 8'h9b, 8'h98, 8'h77, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h74, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h92, 8'h80, 8'h71, 8'h63, 8'h6b, 8'h84, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h66, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h7a, 8'h95, 8'h8f, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h76, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h93, 8'h8d, 8'h8e, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h6d, 8'h36, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h5e, 8'h8b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h65, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h55, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h84, 8'h6d, 8'h5f, 8'h6e, 8'h81, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h64, 8'hc, 8'h0, 8'h16, 8'h76, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h75, 8'h14, 8'h0, 8'h0, 8'h38, 8'h71, 8'h8c, 8'h64, 8'h22, 8'h1, 8'h30, 8'h82, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h71, 8'h5d, 8'h1b, 8'h0, 8'h4d, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h52, 8'he, 8'h22, 8'h75, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h56, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h8c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h72, 8'h2c, 8'h0, 8'h0, 8'h57, 8'h8f, 8'h8d, 8'h5b, 8'h0, 8'h11, 8'h57, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h7c, 8'h73, 8'h85, 8'h9b, 8'h97, 8'h78, 8'h16, 8'h0, 8'h0, 8'h3, 8'h0, 8'h0, 8'h26, 8'h79, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8f, 8'h74, 8'h56, 8'h57, 8'h80, 8'h96, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h36, 8'h76, 8'h50, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h64, 8'h8d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h80, 8'h58, 8'h3b, 8'h3e, 8'h61, 8'h87, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h97, 8'h97, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h84, 8'h66, 8'h3f, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h87, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h65, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h7f, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h76, 8'h4f, 8'h5b, 8'h7b, 8'h95, 8'h9a, 8'h96, 8'h70, 8'h19, 8'h0, 8'h1, 8'h7a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7a, 8'h32, 8'h0, 8'h0, 8'h1a, 8'h55, 8'h14, 8'h0, 8'h2f, 8'h8e, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h63, 8'h2a, 8'h4d, 8'h22, 8'h0, 8'h0, 8'h6b, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h8a, 8'h8c, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h72, 8'h2, 8'h0, 8'h0, 8'h4d, 8'h91, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h60, 8'h8e, 8'h9a, 8'h9a, 8'h8c, 8'h4b, 8'h0, 8'h12, 8'h66, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h75, 8'h6, 8'h0, 8'h1e, 8'h94, 8'h95, 8'h70, 8'h8, 8'h0, 8'h0, 8'h27, 8'h66, 8'h80, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h66, 8'h4b, 8'h61, 8'h88, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h4e, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h54, 8'h87, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h85, 8'h53, 8'hc, 8'h0, 8'h0, 8'h18, 8'h6c, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h74, 8'h72, 8'h83, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8b, 8'h7e, 8'h6a, 8'h50, 8'h28, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h65, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h84, 8'h62, 8'h52, 8'h6e, 8'h9a, 8'h7c, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h58, 8'h13, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h85, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h58, 8'h0, 8'ha, 8'h53, 8'h3a, 8'h0, 8'h0, 8'h4a, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'h30, 8'h0, 8'h0, 8'h26, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h4e, 8'h0, 8'h0, 8'h1c, 8'h5f, 8'h8e, 8'h99, 8'h9b, 8'h9a, 8'h97, 8'h7e, 8'h39, 8'h6, 8'h1b, 8'h7b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h84, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h7, 8'h25, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h47, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h81, 8'h63, 8'h64, 8'h77, 8'h88, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h50, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h66, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h7f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h69, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h45, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h5c, 8'h20, 8'h1c, 8'h4b, 8'h7f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h93, 8'h8e, 8'h8a, 8'h89, 8'h89, 8'h86, 8'h87, 8'h87, 8'h88, 8'h8a, 8'h8d, 8'h90, 8'h89, 8'h74, 8'h44, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h65, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h76, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h88, 8'h79, 8'h60, 8'h49, 8'h24, 8'h0, 8'h0, 8'h24, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8a, 8'h6f, 8'h4f, 8'h3d, 8'h4b, 8'h74, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8d, 8'h4f, 8'h0, 8'h0, 8'h51, 8'h84, 8'h72, 8'h22, 8'h0, 8'h0, 8'h50, 8'h8f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7c, 8'h38, 8'h0, 8'h0, 8'h1e, 8'h73, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h77, 8'h3b, 8'h0, 8'h0, 8'h24, 8'h6d, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h6e, 8'h25, 8'h0, 8'h2a, 8'h7e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h76, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h98, 8'h9b, 8'h9a, 8'h98, 8'h88, 8'h6d, 8'h5e, 8'h68, 8'h7f, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h71, 8'h5d, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h36, 8'h74, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h49, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h79, 8'h1f, 8'h0, 8'h0, 8'h9, 8'h5d, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8f, 8'h7c, 8'h58, 8'h34, 8'h1c, 8'h13, 8'hf, 8'hc, 8'ha, 8'ha, 8'h12, 8'h27, 8'h4b, 8'h71, 8'h8a, 8'h8f, 8'h79, 8'h4f, 8'h9, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h6a, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h67, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h92, 8'h70, 8'h2a, 8'h0, 8'h0, 8'h14, 8'h6a, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h97, 8'h8f, 8'h87, 8'h8b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h4f, 8'ha, 8'h0, 8'h48, 8'h86, 8'h98, 8'h92, 8'h6b, 8'h14, 8'h0, 8'h0, 8'h28, 8'h49, 8'h8a, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7b, 8'h39, 8'h0, 8'h0, 8'h13, 8'h68, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h75, 8'h33, 8'h0, 8'h0, 8'h26, 8'h69, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8e, 8'h5b, 8'hc, 8'h0, 8'h43, 8'h81, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h79, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h5b, 8'h40, 8'h0, 8'h0, 8'ha, 8'h6b, 8'h96, 8'h98, 8'h85, 8'h68, 8'h53, 8'h61, 8'h87, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h7c, 8'h7e, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h70, 8'h8f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h83, 8'h37, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h43, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h8f, 8'h6f, 8'h4d, 8'h2b, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h4f, 8'h78, 8'h8c, 8'h80, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h73, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h76, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h64, 8'ha, 8'h0, 8'h0, 8'h41, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h5a, 8'ha, 8'h0, 8'h40, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h92, 8'h70, 8'h17, 8'h0, 8'h0, 8'h0, 8'h7f, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h82, 8'h3e, 8'h0, 8'h0, 8'h7, 8'h66, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7a, 8'h2d, 8'h0, 8'h0, 8'h42, 8'h7b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h54, 8'h0, 8'h0, 8'h48, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h45, 8'h0, 8'h0, 8'h2b, 8'h74, 8'h57, 8'h62, 8'h7f, 8'h93, 8'h7f, 8'h1c, 8'h0, 8'h0, 8'h12, 8'h84, 8'h85, 8'h63, 8'h53, 8'h6e, 8'h8f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h7e, 8'h91, 8'h7c, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h6d, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7d, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h8f, 8'h6a, 8'h29, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h7a, 8'h8e, 8'h80, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h7f, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h88, 8'h2b, 8'h0, 8'h0, 8'h29, 8'h49, 8'h69, 8'h8c, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h74, 8'h7, 8'h0, 8'h3f, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h72, 8'hf, 8'h0, 8'h2, 8'h87, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h53, 8'h0, 8'h0, 8'h7, 8'h77, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h1d, 8'h0, 8'h0, 8'h4d, 8'h86, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8d, 8'h58, 8'h0, 8'h0, 8'h4a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h72, 8'h0, 8'h0, 8'h1a, 8'h99, 8'h90, 8'h92, 8'h98, 8'h9b, 8'h96, 8'h6c, 8'h3, 8'h0, 8'h0, 8'h43, 8'h48, 8'h63, 8'h84, 8'h92, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h7b, 8'h98, 8'h92, 8'h72, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h5f, 8'h8a, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7d, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h50, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h33, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h99, 8'h8f, 8'h67, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h6c, 8'h88, 8'h71, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h82, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h7a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h1c, 8'h0, 8'h0, 8'h6d, 8'h82, 8'h65, 8'h54, 8'h7b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h4c, 8'h0, 8'h3c, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h7c, 8'h1a, 8'h0, 8'h3a, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h77, 8'h0, 8'h0, 8'ha, 8'h6d, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h74, 8'h16, 8'h0, 8'h0, 8'h3f, 8'h86, 8'h99, 8'h9a, 8'h99, 8'h8c, 8'h64, 8'h27, 8'h50, 8'h83, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h86, 8'h36, 8'h0, 8'h0, 8'h57, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h3b, 8'h2e, 8'h57, 8'h8b, 8'h99, 8'h74, 8'h0, 8'h0, 8'he, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h62, 8'h2b, 8'h14, 8'h3f, 8'h6a, 8'h87, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h8f, 8'h5b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4, 8'h79, 8'h97, 8'h98, 8'h8b, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h81, 8'h95, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7b, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h43, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h43, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h6d, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h62, 8'h7d, 8'h68, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h63, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h73, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6b, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h66, 8'h42, 8'h5f, 8'h8e, 8'h98, 8'h85, 8'h68, 8'h54, 8'h67, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h55, 8'h0, 8'h5, 8'h60, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h80, 8'h2c, 8'h8, 8'h30, 8'h7c, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h79, 8'h2a, 8'h0, 8'h0, 8'h3d, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h76, 8'h2c, 8'h0, 8'h0, 8'h3c, 8'h7b, 8'h99, 8'h9b, 8'h9a, 8'h8b, 8'h5a, 8'h5, 8'h0, 8'h7, 8'h5c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h73, 8'h21, 8'h0, 8'h8, 8'h60, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h72, 8'h0, 8'h0, 8'h0, 8'h24, 8'h2f, 8'h1b, 8'h0, 8'h0, 8'h19, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h75, 8'h51, 8'h44, 8'h68, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h73, 8'h96, 8'h95, 8'h81, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h7a, 8'h93, 8'h99, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h78, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h84, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h84, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h62, 8'h7d, 8'h62, 8'h6, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h71, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h8b, 8'h96, 8'h9a, 8'h9a, 8'h97, 8'h88, 8'h67, 8'h5d, 8'h67, 8'h82, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h49, 8'h0, 8'h0, 8'h2b, 8'h6a, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h79, 8'h31, 8'h9, 8'h2f, 8'h6f, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7c, 8'h3d, 8'h0, 8'h0, 8'h26, 8'h72, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h40, 8'h0, 8'h0, 8'h3c, 8'h7c, 8'h98, 8'h9b, 8'h98, 8'h85, 8'h58, 8'ha, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h60, 8'h14, 8'h0, 8'hd, 8'h61, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h77, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h47, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h7c, 8'h61, 8'h56, 8'h6c, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h69, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6b, 8'h8e, 8'h81, 8'h52, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h92, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h77, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h82, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h85, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h7f, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h70, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h71, 8'h80, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5c, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h80, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h74, 8'h5f, 8'h67, 8'h85, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h66, 8'h10, 8'h0, 8'h0, 8'h20, 8'h5a, 8'h7b, 8'h94, 8'h96, 8'h77, 8'h36, 8'h0, 8'h2b, 8'h6e, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h50, 8'h0, 8'h0, 8'h1c, 8'h6c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h5e, 8'hb, 8'h0, 8'h17, 8'h74, 8'h98, 8'h9b, 8'h9a, 8'h8c, 8'h50, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h58, 8'h3, 8'h0, 8'h12, 8'h65, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h5e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h38, 8'h75, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h83, 8'h56, 8'h64, 8'h80, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h71, 8'h48, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h77, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h78, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h82, 8'h68, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h73, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h84, 8'h66, 8'h56, 8'h80, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h95, 8'h88, 8'h6f, 8'h27, 8'h0, 8'h0, 8'h2c, 8'h78, 8'h7d, 8'h35, 8'h0, 8'h1e, 8'h74, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h77, 8'h19, 8'h0, 8'h4, 8'h74, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7b, 8'h19, 8'h0, 8'h0, 8'h74, 8'h93, 8'h9b, 8'h9a, 8'h94, 8'h64, 8'h0, 8'h0, 8'h0, 8'h35, 8'h6d, 8'h5b, 8'h13, 8'h10, 8'h86, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h4e, 8'h0, 8'h0, 8'h1e, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h89, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h6d, 8'h4f, 8'h75, 8'h8b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h71, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h77, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h73, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h6f, 8'h92, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h98, 8'h7c, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h36, 8'h48, 8'h51, 8'h55, 8'h55, 8'h4c, 8'h34, 8'h6, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h72, 8'h81, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h6e, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8b, 8'h71, 8'h4e, 8'h65, 8'h88, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7e, 8'h5e, 8'h21, 8'h0, 8'h1a, 8'h13, 8'h0, 8'hb, 8'h79, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h1d, 8'h0, 8'h0, 8'h6c, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h2e, 8'h0, 8'h0, 8'h56, 8'h92, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'h1, 8'h0, 8'h0, 8'h30, 8'h7a, 8'h90, 8'h6f, 8'h17, 8'h0, 8'h6a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h84, 8'h43, 8'h0, 8'h0, 8'h21, 8'h6e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h70, 8'h16, 8'h0, 8'h0, 8'h2e, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7d, 8'h63, 8'h5e, 8'h75, 8'h91, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h78, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h7d, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h67, 8'h8f, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h94, 8'h64, 8'h6, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h66, 8'h83, 8'h8c, 8'h8f, 8'h90, 8'h90, 8'h8b, 8'h80, 8'h5a, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5c, 8'h8a, 8'h78, 8'h32, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h6f, 8'h5a, 8'h60, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h6a, 8'h28, 8'h0, 8'h0, 8'h0, 8'h35, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h82, 8'h26, 8'h0, 8'h0, 8'h43, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h57, 8'h0, 8'h0, 8'h40, 8'h8d, 8'h9a, 8'h9b, 8'h9a, 8'h91, 8'h56, 8'h0, 8'h0, 8'h0, 8'h59, 8'h98, 8'h88, 8'h40, 8'hb, 8'h20, 8'h7a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h83, 8'h32, 8'h0, 8'h0, 8'h29, 8'h83, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h54, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h7e, 8'h9b, 8'h94, 8'h75, 8'h5f, 8'h5d, 8'h73, 8'h96, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h79, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h62, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h76, 8'h23, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h62, 8'h8d, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h91, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h64, 8'h8c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h59, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h40, 8'h82, 8'h8c, 8'h6e, 8'h3b, 8'h21, 8'h2f, 8'h66, 8'h93, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h85, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h90, 8'h72, 8'h5f, 8'h60, 8'h7b, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h92, 8'h70, 8'h26, 8'h0, 8'h1a, 8'h6a, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h51, 8'h0, 8'h0, 8'h34, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h63, 8'h11, 8'h0, 8'h33, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h62, 8'h0, 8'h0, 8'h0, 8'h44, 8'h7c, 8'h52, 8'h7, 8'h16, 8'h63, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h80, 8'h31, 8'h0, 8'h0, 8'h4a, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h47, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h8a, 8'h78, 8'h5a, 8'h5d, 8'h78, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h96, 8'h72, 8'h16, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h5e, 8'h8c, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h98, 8'h8c, 8'h49, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h55, 8'h86, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h82, 8'h52, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h62, 8'h8c, 8'h8c, 8'h7e, 8'h75, 8'h7e, 8'h8e, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h7a, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h79, 8'h61, 8'h5a, 8'h81, 8'h93, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h7a, 8'h4e, 8'h5c, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h63, 8'hc, 8'h0, 8'h26, 8'h74, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h6d, 8'h22, 8'h0, 8'h16, 8'h68, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h47, 8'h0, 8'h0, 8'h0, 8'h23, 8'h0, 8'h0, 8'h49, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h80, 8'h2c, 8'h0, 8'h0, 8'h5a, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h86, 8'h48, 8'h0, 8'h0, 8'h14, 8'h56, 8'h46, 8'h66, 8'h86, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h76, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'hf, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h55, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h96, 8'h6e, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h5f, 8'h8c, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h7e, 8'h32, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h32, 8'h7d, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h7f, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h82, 8'h98, 8'h97, 8'h95, 8'h97, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h7d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h8c, 8'h70, 8'h4f, 8'h79, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h92, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h76, 8'h25, 8'h0, 8'h0, 8'h5d, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h74, 8'h29, 8'h0, 8'h1, 8'h61, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h86, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h89, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h73, 8'h22, 8'h0, 8'h0, 8'h55, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h83, 8'h39, 8'h0, 8'h0, 8'h38, 8'h7a, 8'h8c, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h79, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h37, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h95, 8'h6c, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h62, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h5c, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5c, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h7c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h76, 8'hf, 8'h0, 8'h0, 8'h55, 8'h89, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h91, 8'h7a, 8'h5b, 8'h6a, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h28, 8'h0, 8'h0, 8'h56, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7c, 8'h2e, 8'h0, 8'h0, 8'h5a, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h54, 8'h2a, 8'h2d, 8'h54, 8'h84, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h6c, 8'h1a, 8'h0, 8'h0, 8'h4c, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h67, 8'h27, 8'h2f, 8'h6d, 8'h94, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7d, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h4c, 8'h69, 8'h79, 8'h6a, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7d, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h95, 8'h6a, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h69, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h7c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h70, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h78, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h77, 8'h61, 8'h75, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h76, 8'h61, 8'h64, 8'h7f, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h3b, 8'h0, 8'h0, 8'h4a, 8'h89, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h36, 8'h0, 8'h0, 8'h4d, 8'h90, 8'h99, 8'h9a, 8'h8f, 8'h83, 8'h8a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8e, 8'h83, 8'h80, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h6a, 8'h15, 8'h0, 8'h0, 8'h3a, 8'h6a, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h7a, 8'h62, 8'h5e, 8'h77, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h80, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h1d, 8'h34, 8'h46, 8'h5b, 8'h72, 8'h86, 8'h91, 8'h95, 8'h8e, 8'h6f, 8'h23, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h99, 8'h9a, 8'h95, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h71, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'h23, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h73, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h77, 8'h5d, 8'h5b, 8'h79, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h56, 8'h0, 8'h0, 8'h26, 8'h8e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h7c, 8'h3f, 8'h0, 8'h0, 8'h47, 8'h92, 8'h9a, 8'h92, 8'h76, 8'h52, 8'h3c, 8'h4e, 8'h7e, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h62, 8'h0, 8'h0, 8'h0, 8'h19, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h75, 8'h58, 8'h5b, 8'h80, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h27, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h5c, 8'h72, 8'h7f, 8'h89, 8'h8f, 8'h95, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h8d, 8'h60, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h85, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h66, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h78, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h74, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h6d, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h66, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h7a, 8'h55, 8'h54, 8'h79, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h6d, 8'hb, 8'h0, 8'h9, 8'h60, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h81, 8'h38, 8'h0, 8'h0, 8'h46, 8'h90, 8'h9b, 8'h97, 8'h70, 8'h10, 8'h0, 8'h0, 8'h0, 8'h44, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h78, 8'h2, 8'h0, 8'h0, 8'h0, 8'h64, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h91, 8'h6c, 8'h4b, 8'h5a, 8'h89, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h36, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4f, 8'h86, 8'h93, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h40, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h36, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h70, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h52, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h7c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h73, 8'h13, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h83, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h87, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h91, 8'h8d, 8'h8e, 8'h94, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h85, 8'h5d, 8'h51, 8'h73, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h3d, 8'h0, 8'h0, 8'h4f, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h35, 8'h0, 8'h0, 8'h42, 8'h84, 8'h9b, 8'h9b, 8'h7d, 8'h9, 8'h0, 8'h0, 8'h16, 8'h0, 8'h7, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7f, 8'h15, 8'h0, 8'h0, 8'h0, 8'h0, 8'h60, 8'h9a, 8'h9a, 8'h9b, 8'h91, 8'h65, 8'h56, 8'h69, 8'h8a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8c, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5c, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h72, 8'h16, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h80, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6e, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h60, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h76, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h76, 8'h42, 8'h27, 8'h34, 8'h55, 8'h75, 8'h86, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h86, 8'h6b, 8'h57, 8'h6b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h4b, 8'h0, 8'h0, 8'h42, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h3b, 8'h0, 8'h0, 8'h3a, 8'h7f, 8'h98, 8'h97, 8'h7e, 8'h2e, 8'h0, 8'h0, 8'h30, 8'h6b, 8'h41, 8'h0, 8'h31, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h73, 8'h19, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h36, 8'h7d, 8'h9b, 8'h9a, 8'h8c, 8'h66, 8'h60, 8'h6f, 8'h8a, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h60, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h50, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h79, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6f, 8'hf, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h81, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h63, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h71, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7e, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h66, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8f, 8'h49, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h88, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h89, 8'h73, 8'h64, 8'h6b, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h51, 8'h0, 8'h0, 8'h25, 8'h79, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h48, 8'h0, 8'h0, 8'h2e, 8'h86, 8'h96, 8'h9a, 8'h8e, 8'h57, 8'h0, 8'h0, 8'h1b, 8'h71, 8'h95, 8'h75, 8'h12, 8'h7, 8'h38, 8'h6f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6d, 8'h20, 8'h0, 8'h0, 8'h3, 8'h54, 8'h8b, 8'h87, 8'h95, 8'h98, 8'h88, 8'h6c, 8'h5d, 8'h74, 8'h8d, 8'h98, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h68, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4a, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h48, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h70, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h80, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h83, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h78, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h88, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5e, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h48, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h38, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h79, 8'h5f, 8'h73, 8'h8b, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h56, 8'h8, 8'h0, 8'h1a, 8'h6f, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h8e, 8'h5d, 8'h0, 8'h0, 8'h2c, 8'h7e, 8'h98, 8'h9b, 8'h96, 8'h75, 8'h24, 8'h0, 8'h0, 8'h4c, 8'h97, 8'h9b, 8'h86, 8'h26, 8'h0, 8'h0, 8'h32, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h70, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h55, 8'h93, 8'h99, 8'h99, 8'h96, 8'h89, 8'h6b, 8'h54, 8'h80, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'hc, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h36, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7b, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h58, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8b, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7f, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h7e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h6e, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h82, 8'h5b, 8'h6f, 8'h89, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h73, 8'hb, 8'h0, 8'h1f, 8'h78, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h5d, 8'h0, 8'h0, 8'h38, 8'h82, 8'h98, 8'h9b, 8'h9b, 8'h8b, 8'h34, 8'h0, 8'h0, 8'h35, 8'h7e, 8'h9b, 8'h9b, 8'h7e, 8'h10, 8'h0, 8'h0, 8'h41, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h14, 8'h0, 8'h0, 8'h0, 8'h53, 8'h91, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h60, 8'h5f, 8'h90, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8b, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h69, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h68, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h6a, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h93, 8'h72, 8'h23, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h77, 8'h27, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h86, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h84, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h7c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h59, 8'h62, 8'h8b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h42, 8'h0, 8'h24, 8'h7a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h51, 8'h0, 8'h0, 8'h2b, 8'h73, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h2a, 8'h0, 8'h0, 8'h3a, 8'h80, 8'h99, 8'h77, 8'h1b, 8'h0, 8'h0, 8'h11, 8'h81, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h84, 8'h1e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h6a, 8'h9b, 8'h96, 8'h80, 8'h5f, 8'h6a, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h7e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h56, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h45, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h32, 8'h75, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h7f, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h41, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h71, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8d, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7f, 8'h62, 8'h5c, 8'h80, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8c, 8'h55, 8'h0, 8'h0, 8'h4a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h53, 8'ha, 8'h0, 8'h25, 8'h6f, 8'h90, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h57, 8'h0, 8'h0, 8'h0, 8'h32, 8'h3d, 8'he, 8'h0, 8'h0, 8'h7, 8'h5f, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h74, 8'h21, 8'h0, 8'h0, 8'h0, 8'h18, 8'h9, 8'h0, 8'h4d, 8'h90, 8'h7a, 8'h60, 8'h6a, 8'h85, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h77, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h7f, 8'h36, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h49, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h32, 8'h6f, 8'h8e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h83, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6a, 8'hc, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5f, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h81, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7e, 8'h60, 8'h5b, 8'h79, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h56, 8'h2, 8'h0, 8'h31, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h65, 8'h11, 8'h0, 8'h1e, 8'h76, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h86, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h58, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h71, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h43, 8'h27, 8'h0, 8'h39, 8'h77, 8'h5e, 8'h63, 8'h87, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h72, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h61, 8'h86, 8'h95, 8'h99, 8'h9a, 8'h98, 8'h92, 8'h7a, 8'h49, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h63, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h64, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h66, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h71, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h80, 8'h5c, 8'h5e, 8'h76, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h61, 8'hf, 8'h0, 8'h25, 8'h76, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h8f, 8'h6b, 8'h1f, 8'h0, 8'h15, 8'h68, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h63, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h77, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h5a, 8'h5f, 8'h8e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h62, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h69, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h8a, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h52, 8'h71, 8'h7c, 8'h80, 8'h7c, 8'h6a, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h7b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h60, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h67, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h86, 8'h5e, 8'h5a, 8'h74, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h75, 8'h1b, 8'h0, 8'h1, 8'h7e, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h93, 8'h60, 8'h0, 8'h0, 8'h4, 8'h55, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h5d, 8'h0, 8'h0, 8'h7, 8'h78, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7f, 8'h18, 8'h0, 8'h0, 8'h0, 8'h49, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h16, 8'h63, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h97, 8'h9b, 8'h9a, 8'h95, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h9, 8'h6, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h16, 8'h6f, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h87, 8'h61, 8'h51, 8'h6b, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h85, 8'h27, 8'h0, 8'h0, 8'h43, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h4d, 8'h0, 8'h0, 8'h1a, 8'h5a, 8'h8a, 8'h9a, 8'h91, 8'h78, 8'h88, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h69, 8'h56, 8'h6c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h81, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h57, 8'h86, 8'h6e, 8'h21, 8'h0, 8'h0, 8'hb, 8'h55, 8'h89, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h98, 8'h97, 8'h97, 8'h96, 8'h96, 8'h95, 8'h95, 8'h94, 8'h93, 8'h93, 8'h93, 8'h92, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h93, 8'h93, 8'h90, 8'h91, 8'h91, 8'h91, 8'h92, 8'h91, 8'h8f, 8'h8e, 8'h8d, 8'h8e, 8'h8e, 8'h90, 8'h91, 8'h91, 8'h92, 8'h91, 8'h8f, 8'h8e, 8'h8e, 8'h8d, 8'h8f, 8'h91, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h93, 8'h92, 8'h93, 8'h95, 8'h96, 8'h96, 8'h95, 8'h95, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h95, 8'h96, 8'h96, 8'h96, 8'h95, 8'h95, 8'h96, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h97, 8'h98, 8'h98, 8'h98, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h74, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h97, 8'h72, 8'h6, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h65, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h78, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h92, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h85, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h98, 8'h98, 8'h98, 8'h97, 8'h96, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h95, 8'h94, 8'h93, 8'h93, 8'h92, 8'h91, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h90, 8'h8e, 8'h8d, 8'h8d, 8'h8e, 8'h8d, 8'h8d, 8'h8e, 8'h8e, 8'h8e, 8'h8c, 8'h8b, 8'h8c, 8'h8c, 8'h8d, 8'h8e, 8'h8c, 8'h8d, 8'h8e, 8'h8e, 8'h8d, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8a, 8'h8a, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8d, 8'h8d, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8b, 8'h8c, 8'h8c, 8'h8c, 8'h8e, 8'h8e, 8'h8e, 8'h8d, 8'h8d, 8'h8f, 8'h91, 8'h92, 8'h91, 8'h94, 8'h95, 8'h96, 8'h96, 8'h96, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h84, 8'h67, 8'h54, 8'h6d, 8'h91, 8'h9b, 8'h99, 8'h8c, 8'h58, 8'h0, 8'h0, 8'h2e, 8'h81, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h52, 8'h7, 8'h0, 8'h28, 8'h67, 8'h89, 8'h84, 8'h5e, 8'h21, 8'h10, 8'h29, 8'h62, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h95, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h79, 8'h29, 8'h0, 8'h0, 8'h0, 8'h52, 8'h8f, 8'h98, 8'h8f, 8'h5a, 8'h12, 8'h11, 8'h54, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h8a, 8'h7c, 8'h72, 8'h6f, 8'h6f, 8'h6d, 8'h6b, 8'h6b, 8'h68, 8'h66, 8'h64, 8'h63, 8'h62, 8'h5d, 8'h5d, 8'h5a, 8'h57, 8'h55, 8'h54, 8'h52, 8'h50, 8'h50, 8'h4f, 8'h4d, 8'h4b, 8'h49, 8'h47, 8'h47, 8'h47, 8'h45, 8'h42, 8'h41, 8'h41, 8'h41, 8'h41, 8'h43, 8'h43, 8'h41, 8'h41, 8'h40, 8'h41, 8'h42, 8'h40, 8'h3b, 8'h37, 8'h36, 8'h37, 8'h39, 8'h3d, 8'h41, 8'h43, 8'h42, 8'h40, 8'h3b, 8'h39, 8'h37, 8'h37, 8'h3a, 8'h41, 8'h46, 8'h47, 8'h47, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h47, 8'h48, 8'h4b, 8'h4e, 8'h4e, 8'h4e, 8'h4e, 8'h4f, 8'h4e, 8'h4d, 8'h4d, 8'h4d, 8'h4e, 8'h4e, 8'h4e, 8'h4d, 8'h4e, 8'h4e, 8'h4e, 8'h4d, 8'h4d, 8'h4e, 8'h50, 8'h52, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h52, 8'h54, 8'h55, 8'h55, 8'h56, 8'h57, 8'h58, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h62, 8'h6b, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8a, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9a, 8'h89, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h79, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h81, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h52, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h52, 8'h90, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h6b, 8'h66, 8'h64, 8'h63, 8'h61, 8'h60, 8'h5e, 8'h5e, 8'h5c, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h58, 8'h56, 8'h55, 8'h55, 8'h53, 8'h50, 8'h50, 8'h50, 8'h4f, 8'h4e, 8'h4e, 8'h4e, 8'h4d, 8'h4b, 8'h49, 8'h47, 8'h46, 8'h44, 8'h42, 8'h41, 8'h42, 8'h42, 8'h42, 8'h42, 8'h41, 8'h3d, 8'h39, 8'h37, 8'h37, 8'h37, 8'h36, 8'h37, 8'h38, 8'h38, 8'h36, 8'h34, 8'h31, 8'h31, 8'h32, 8'h35, 8'h36, 8'h36, 8'h36, 8'h37, 8'h37, 8'h34, 8'h31, 8'h30, 8'h30, 8'h30, 8'h2f, 8'h2f, 8'h30, 8'h30, 8'h2f, 8'h2f, 8'h2f, 8'h30, 8'h32, 8'h32, 8'h30, 8'h2f, 8'h2f, 8'h2f, 8'h30, 8'h30, 8'h2f, 8'h2f, 8'h2f, 8'h30, 8'h30, 8'h2f, 8'h2f, 8'h30, 8'h31, 8'h33, 8'h34, 8'h38, 8'h37, 8'h37, 8'h37, 8'h37, 8'h3c, 8'h42, 8'h44, 8'h44, 8'h47, 8'h4b, 8'h4e, 8'h4f, 8'h51, 8'h54, 8'h5a, 8'h5d, 8'h60, 8'h62, 8'h65, 8'h6a, 8'h79, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h84, 8'h67, 8'h54, 8'h6d, 8'h8a, 8'h99, 8'h6e, 8'h9, 8'h0, 8'h1c, 8'h6f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8f, 8'h5d, 8'hc, 8'h0, 8'h26, 8'h7c, 8'h94, 8'h8f, 8'h5c, 8'h5, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h6d, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h71, 8'h28, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h93, 8'h9a, 8'h98, 8'h88, 8'h67, 8'h4b, 8'h61, 8'h88, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h68, 8'h40, 8'h23, 8'h16, 8'h14, 8'h10, 8'h7, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h81, 8'h43, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h96, 8'h9b, 8'h94, 8'h72, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4, 8'h5a, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h45, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h57, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h52, 8'h90, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h61, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h93, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h5c, 8'h4, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h85, 8'h62, 8'h56, 8'h6e, 8'h76, 8'h41, 8'h0, 8'h0, 8'h56, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8f, 8'h64, 8'h8, 8'h0, 8'h21, 8'h72, 8'h99, 8'h9a, 8'h88, 8'h25, 8'h0, 8'h0, 8'h38, 8'h1b, 8'h0, 8'h19, 8'h80, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h73, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h52, 8'h91, 8'h9b, 8'h9a, 8'h8c, 8'h6b, 8'h53, 8'h62, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h85, 8'h7e, 8'h7d, 8'h7b, 8'h73, 8'h70, 8'h66, 8'h5c, 8'h52, 8'h47, 8'h36, 8'h22, 8'hd, 8'h4, 8'h1, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2, 8'h3, 8'h2, 8'h4, 8'h5, 8'h7, 8'h7, 8'h16, 8'h3c, 8'h69, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h65, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h71, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h72, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h72, 8'h9b, 8'h99, 8'h90, 8'h64, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h7c, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h8f, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h69, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h74, 8'h5d, 8'h52, 8'h45, 8'h3d, 8'h33, 8'h25, 8'h16, 8'h7, 8'h3, 8'h5, 8'h3, 8'h2, 8'h3, 8'h3, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h6, 8'h19, 8'h36, 8'h44, 8'h53, 8'h6d, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h67, 8'h50, 8'h3c, 8'hd, 8'h0, 8'h40, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5b, 8'h0, 8'h0, 8'h1d, 8'h69, 8'h95, 8'h9b, 8'h9a, 8'h7f, 8'h18, 8'h0, 8'h0, 8'h6f, 8'h76, 8'h2a, 8'h0, 8'hc, 8'h7c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h80, 8'h11, 8'h0, 8'h0, 8'h0, 8'h63, 8'h8f, 8'h9a, 8'h9b, 8'h8f, 8'h63, 8'h52, 8'h69, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h76, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h60, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h57, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8c, 8'h9b, 8'h9a, 8'h99, 8'h8e, 8'h64, 8'h23, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h70, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h67, 8'he, 8'h0, 8'h0, 8'h0, 8'h14, 8'h67, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6c, 8'h16, 8'h0, 8'h0, 8'h0, 8'h3, 8'h62, 8'h93, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h98, 8'h98, 8'h99, 8'h99, 8'h99, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h99, 8'h98, 8'h98, 8'h98, 8'h99, 8'h99, 8'h99, 8'h98, 8'h98, 8'h98, 8'h99, 8'h99, 8'h98, 8'h98, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h63, 8'h22, 8'h0, 8'h1, 8'h6e, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h58, 8'h9, 8'h0, 8'h1b, 8'h63, 8'h8e, 8'h9b, 8'h9b, 8'h8a, 8'h40, 8'h0, 8'h0, 8'h25, 8'h84, 8'h94, 8'h6d, 8'h1e, 8'h0, 8'h10, 8'h6a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7a, 8'h14, 8'h0, 8'h0, 8'h6, 8'h64, 8'h8e, 8'h9b, 8'h99, 8'h8b, 8'h67, 8'h55, 8'h6b, 8'h89, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7e, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h73, 8'h45, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h71, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h7e, 8'h46, 8'h1f, 8'h23, 8'h38, 8'h5d, 8'h85, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h81, 8'h42, 8'h0, 8'h0, 8'h0, 8'h41, 8'h7d, 8'h95, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h62, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h65, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h5e, 8'h2c, 8'h32, 8'h80, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h5f, 8'h13, 8'h0, 8'h1a, 8'h64, 8'h8c, 8'h9a, 8'h9b, 8'h9a, 8'h7c, 8'ha, 8'h0, 8'h0, 8'h69, 8'h92, 8'h9a, 8'h8c, 8'h40, 8'h0, 8'h0, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h70, 8'h1c, 8'h0, 8'h0, 8'hb, 8'h5d, 8'h95, 8'h9b, 8'h97, 8'h88, 8'h6a, 8'h54, 8'h6c, 8'h89, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h45, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h6b, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h7e, 8'h5f, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h36, 8'h6c, 8'h8e, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h77, 8'h67, 8'h6d, 8'h7a, 8'h88, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h70, 8'h3e, 8'h25, 8'h43, 8'h73, 8'h90, 8'h9a, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h64, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h50, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h86, 8'h69, 8'h50, 8'h6c, 8'h8b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h77, 8'h1f, 8'h0, 8'h14, 8'h6b, 8'h90, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h76, 8'h0, 8'h0, 8'h0, 8'h63, 8'h8e, 8'h92, 8'h6f, 8'h1c, 8'h0, 8'h0, 8'h5c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h71, 8'h21, 8'h0, 8'h0, 8'h9, 8'h5a, 8'h94, 8'h9b, 8'h98, 8'h8a, 8'h6d, 8'h55, 8'h67, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h87, 8'h58, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h8a, 8'h71, 8'h3f, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h30, 8'h4c, 8'h60, 8'h78, 8'h8e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h92, 8'h8f, 8'h92, 8'h96, 8'h98, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h7a, 8'h71, 8'h7f, 8'h91, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h99, 8'h98, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h76, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h60, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h8b, 8'h69, 8'h58, 8'h70, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h49, 8'h0, 8'hb, 8'h5b, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h19, 8'h0, 8'h0, 8'h0, 8'h64, 8'h6a, 8'h1b, 8'h0, 8'h0, 8'h39, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h7a, 8'h20, 8'h0, 8'h0, 8'h0, 8'h5e, 8'h94, 8'h9b, 8'h9b, 8'h8c, 8'h6b, 8'h53, 8'h62, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h84, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h86, 8'h66, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h91, 8'h7a, 8'h59, 8'h3f, 8'h30, 8'h27, 8'h1b, 8'h13, 8'he, 8'h14, 8'h1f, 8'h2e, 8'h41, 8'h61, 8'h7c, 8'h8b, 8'h91, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h95, 8'h97, 8'h9a, 8'h9b, 8'h98, 8'h97, 8'h98, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h6f, 8'h59, 8'h3d, 8'h2e, 8'h31, 8'h4b, 8'h5f, 8'h83, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8e, 8'h69, 8'h59, 8'h6d, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h8f, 8'h58, 8'h0, 8'h0, 8'h47, 8'h8e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h71, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h73, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h84, 8'h22, 8'h0, 8'h0, 8'h0, 8'h65, 8'h91, 8'h9a, 8'h9b, 8'h91, 8'h67, 8'h55, 8'h69, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h38, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h91, 8'h7c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h42, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h8a, 8'h82, 8'h7c, 8'h78, 8'h70, 8'h69, 8'h65, 8'h69, 8'h70, 8'h7a, 8'h83, 8'h8e, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h8b, 8'h8e, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h6b, 8'h56, 8'h64, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h59, 8'h0, 8'h0, 8'h3c, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h6a, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h67, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7e, 8'h22, 8'h0, 8'h0, 8'h0, 8'h61, 8'h8f, 8'h99, 8'h99, 8'h8d, 8'h6d, 8'h54, 8'h6b, 8'h8a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h66, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h43, 8'h89, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h83, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h98, 8'h97, 8'h96, 8'h94, 8'h90, 8'h90, 8'h91, 8'h94, 8'h95, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h87, 8'h67, 8'h51, 8'h6c, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h60, 8'he, 8'h0, 8'h25, 8'h78, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h6d, 8'h27, 8'h0, 8'h0, 8'h1f, 8'h5c, 8'h94, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7d, 8'h37, 8'h0, 8'h0, 8'h0, 8'h50, 8'h95, 8'h9a, 8'h99, 8'h8b, 8'h6f, 8'h56, 8'h68, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h51, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h58, 8'h57, 8'h86, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h84, 8'h63, 8'h52, 8'h71, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7a, 8'h47, 8'h4a, 8'h7b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h68, 8'h17, 8'h0, 8'h12, 8'h75, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h84, 8'h65, 8'h61, 8'h78, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h47, 8'h0, 8'h0, 8'h0, 8'h51, 8'h94, 8'h9a, 8'h9a, 8'h8e, 8'h73, 8'h5a, 8'h63, 8'h8b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h61, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h70, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h85, 8'h5d, 8'h58, 8'h74, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h76, 8'h2f, 8'h0, 8'h0, 8'h50, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'h13, 8'h0, 8'h13, 8'h74, 8'h95, 8'h9a, 8'h9b, 8'h98, 8'h93, 8'h90, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h95, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h5c, 8'h5, 8'h0, 8'h0, 8'h54, 8'h92, 8'h9b, 8'h9b, 8'h93, 8'h77, 8'h59, 8'h5f, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h6c, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h36, 8'h6e, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h89, 8'h5f, 8'h58, 8'h73, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h82, 8'h29, 8'h0, 8'h0, 8'h0, 8'h34, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'h2e, 8'h0, 8'h15, 8'h64, 8'h95, 8'h9a, 8'h9b, 8'h97, 8'h7e, 8'h45, 8'h23, 8'h6b, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6a, 8'h10, 8'h0, 8'h0, 8'h4c, 8'h88, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h5b, 8'h64, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h81, 8'h68, 8'h54, 8'h43, 8'h39, 8'h3b, 8'h4b, 8'h69, 8'h89, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h86, 8'h62, 8'h58, 8'h76, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h78, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h7f, 8'h76, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h52, 8'h0, 8'h6, 8'h51, 8'h8d, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h49, 8'h0, 8'h0, 8'hc, 8'h58, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h93, 8'h6d, 8'h14, 8'h0, 8'h0, 8'h38, 8'h84, 8'h97, 8'h99, 8'h96, 8'h85, 8'h5e, 8'h6a, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h96, 8'h90, 8'h8a, 8'h89, 8'h90, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h83, 8'h62, 8'h57, 8'h7d, 8'h94, 8'h9b, 8'h99, 8'h8a, 8'h42, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h0, 8'h21, 8'h72, 8'h9b, 8'h94, 8'h70, 8'h45, 8'h24, 8'h11, 8'h3, 8'he, 8'h5e, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8e, 8'h5d, 8'he, 8'h0, 8'h41, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h5e, 8'he, 8'h0, 8'h4, 8'h0, 8'hf, 8'h4d, 8'h7b, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h6d, 8'h1b, 8'h0, 8'h0, 8'h33, 8'h7f, 8'h96, 8'h9a, 8'h94, 8'h7f, 8'h65, 8'h67, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h80, 8'h5f, 8'h60, 8'h82, 8'h94, 8'h89, 8'h55, 8'h0, 8'h0, 8'h0, 8'h34, 8'h60, 8'h0, 8'h0, 8'h32, 8'h4d, 8'h3b, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h47, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h67, 8'h18, 8'h0, 8'h21, 8'h78, 8'h98, 8'h9a, 8'h9b, 8'h98, 8'h81, 8'h2b, 8'h0, 8'hb, 8'h68, 8'h29, 8'h0, 8'h0, 8'h37, 8'h79, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h6e, 8'h20, 8'h0, 8'h0, 8'h33, 8'h83, 8'h98, 8'h9a, 8'h96, 8'h81, 8'h64, 8'h5b, 8'h8b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h82, 8'h5a, 8'h6b, 8'h7f, 8'h63, 8'h8, 8'h0, 8'h0, 8'h2e, 8'h7d, 8'h7b, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h80, 8'h1b, 8'h0, 8'h18, 8'h84, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h64, 8'h9, 8'h0, 8'h4d, 8'h8d, 8'h7c, 8'h1c, 8'h0, 8'h0, 8'h50, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h78, 8'h24, 8'h0, 8'h0, 8'h33, 8'h7b, 8'h99, 8'h9b, 8'h9a, 8'h8c, 8'h65, 8'h5d, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h59, 8'h58, 8'h2c, 8'h0, 8'h0, 8'h32, 8'h7c, 8'h98, 8'h93, 8'h64, 8'hb, 8'h0, 8'h0, 8'h11, 8'h5e, 8'h75, 8'h45, 8'h0, 8'h0, 8'h18, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h47, 8'h0, 8'h15, 8'h77, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h73, 8'h9, 8'h0, 8'h19, 8'h88, 8'h98, 8'h87, 8'h26, 8'h0, 8'h0, 8'h73, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h27, 8'h0, 8'h0, 8'h39, 8'h78, 8'h95, 8'h9b, 8'h9b, 8'h90, 8'h66, 8'h68, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7f, 8'h50, 8'h3, 8'h0, 8'h18, 8'h6c, 8'h96, 8'h9b, 8'h9a, 8'h8f, 8'h75, 8'h67, 8'h6a, 8'h78, 8'h90, 8'h88, 8'h34, 8'h0, 8'h0, 8'h55, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h74, 8'h3, 8'h0, 8'h41, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h75, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h8c, 8'h6e, 8'h14, 8'h0, 8'h3b, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h2f, 8'h0, 8'h0, 8'h17, 8'h76, 8'h93, 8'h9b, 8'h9a, 8'h8d, 8'h66, 8'h69, 8'h83, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h70, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h13, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h58, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h70, 8'h6f, 8'h71, 8'h70, 8'h3f, 8'h3f, 8'h71, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h75, 8'h38, 8'he, 8'h63, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h97, 8'h97, 8'h98, 8'h98, 8'h99, 8'h83, 8'h22, 8'h0, 8'h0, 8'h6b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h71, 8'h0, 8'h0, 8'h37, 8'h8b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h88, 8'h40, 8'h16, 8'h0, 8'h0, 8'h40, 8'h22, 8'h0, 8'h9, 8'h7a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8b, 8'h50, 8'h0, 8'h0, 8'h3, 8'h62, 8'h92, 8'h9a, 8'h98, 8'h8b, 8'h6c, 8'h5b, 8'h7e, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h70, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h31, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h86, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h4b, 8'h9b, 8'h9b, 8'h9b, 8'h6f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h74, 8'h4f, 8'h70, 8'h8e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h72, 8'h13, 8'h0, 8'h3, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h2a, 8'h0, 8'h7, 8'h57, 8'h8b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h80, 8'h43, 8'h0, 8'h0, 8'h0, 8'h0, 8'h33, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h68, 8'h0, 8'h0, 8'h0, 8'h47, 8'h95, 8'h99, 8'h99, 8'h8d, 8'h6c, 8'h54, 8'h79, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h70, 8'h71, 8'h70, 8'h70, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h22, 8'h0, 8'h0, 8'h2, 8'h4b, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h2, 8'h13, 8'h0, 8'h0, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h0, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h71, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h0, 8'h0, 8'h3f, 8'h3f, 8'h4d, 8'h70, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h70, 8'h70, 8'h70, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7c, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h74, 8'h56, 8'h76, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h66, 8'ha, 8'h0, 8'h22, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h91, 8'h80, 8'h7e, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7b, 8'h22, 8'h0, 8'h0, 8'h5c, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h88, 8'h4b, 8'h0, 8'h0, 8'h27, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7e, 8'h34, 8'h0, 8'h0, 8'h3a, 8'h90, 8'h9b, 8'h9b, 8'h92, 8'h6b, 8'h56, 8'h70, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2, 8'h0, 8'h0, 8'h0, 8'h2, 8'h31, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h13, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2, 8'h4c, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h6f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h70, 8'h2, 8'h0, 8'h0, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h57, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h0, 8'h0, 8'h1, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h0, 8'h22, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h3e, 8'h0, 8'h0, 8'h13, 8'h9b, 8'h71, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h71, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h6a, 8'h54, 8'h72, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h71, 8'h13, 8'h0, 8'h4, 8'h74, 8'h97, 8'h98, 8'h98, 8'h92, 8'h65, 8'h17, 8'h11, 8'h67, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6f, 8'h22, 8'h0, 8'h0, 8'h2f, 8'h76, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h5f, 8'h5c, 8'h7a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h78, 8'h2e, 8'h0, 8'h0, 8'h2e, 8'h7b, 8'h9b, 8'h9a, 8'h94, 8'h71, 8'h59, 8'h66, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2, 8'h0, 8'h23, 8'h12, 8'h0, 8'h0, 8'h0, 8'h7b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h2, 8'h3f, 8'h2, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h70, 8'h0, 8'h0, 8'h70, 8'h71, 8'h70, 8'h70, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h4c, 8'h0, 8'h0, 8'h13, 8'h4c, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h0, 8'h31, 8'h64, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h0, 8'h0, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9a, 8'h23, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h64, 8'h0, 8'h0, 8'h71, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h0, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h3, 8'h1, 8'h3f, 8'h3f, 8'h0, 8'h0, 8'h22, 8'h40, 8'h13, 8'h1, 8'h3, 8'h9b, 8'h9b, 8'h7a, 8'h0, 8'h0, 8'h3, 8'h58, 8'h70, 8'h71, 8'h30, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h0, 8'h31, 8'h6f, 8'h9b, 8'h7a, 8'h3, 8'h2, 8'h23, 8'h3f, 8'h1, 8'h0, 8'h2, 8'h3f, 8'h22, 8'h2, 8'h2, 8'h58, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h71, 8'h0, 8'h0, 8'h3f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h71, 8'h0, 8'h0, 8'h40, 8'h22, 8'h0, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h58, 8'h2, 8'h2, 8'h31, 8'h3f, 8'h1, 8'h0, 8'h2, 8'h40, 8'h21, 8'h2, 8'h2, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h66, 8'h5b, 8'h74, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h81, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h38, 8'h0, 8'h0, 8'h8, 8'h7a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h6b, 8'h24, 8'h0, 8'h0, 8'h13, 8'h5b, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h97, 8'h94, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h82, 8'h31, 8'h0, 8'h0, 8'h21, 8'h72, 8'h94, 8'h9a, 8'h95, 8'h7a, 8'h5b, 8'h65, 8'h85, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h91, 8'h13, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9b, 8'h71, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h65, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3, 8'h0, 8'h22, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h40, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h3, 8'h9b, 8'h3e, 8'h0, 8'h1, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h0, 8'h0, 8'h32, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h0, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h31, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h86, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h13, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h80, 8'h61, 8'h5a, 8'h7f, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h53, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h74, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h71, 8'h26, 8'h0, 8'h0, 8'h0, 8'h58, 8'h8a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h42, 8'h0, 8'h0, 8'h1a, 8'h72, 8'h91, 8'h9a, 8'h97, 8'h84, 8'h5e, 8'h63, 8'h7f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h86, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h9a, 8'h3f, 8'h0, 8'h40, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h1, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h13, 8'h0, 8'h13, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h31, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h13, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h57, 8'h0, 8'h22, 8'h3f, 8'h0, 8'h2, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h59, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h7a, 8'h5c, 8'h5b, 8'h88, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h82, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h77, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7d, 8'h28, 8'h0, 8'h0, 8'h0, 8'h53, 8'h7d, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h5e, 8'h0, 8'h0, 8'hf, 8'h77, 8'h95, 8'h9a, 8'h99, 8'h8c, 8'h6e, 8'h59, 8'h82, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h71, 8'h9a, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h13, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h57, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h3, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h0, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h86, 8'h91, 8'h0, 8'h0, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h77, 8'h50, 8'h71, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h16, 8'h0, 8'h1d, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h44, 8'h0, 8'h0, 8'h0, 8'h20, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h60, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h97, 8'h9b, 8'h9b, 8'h94, 8'h71, 8'h4f, 8'h89, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3, 8'h0, 8'h6e, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h40, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h40, 8'h9a, 8'h4c, 8'h0, 8'h0, 8'h7c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h2, 8'h2, 8'h3, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h3, 8'h0, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h0, 8'h0, 8'h0, 8'h22, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h3f, 8'h86, 8'h21, 8'h0, 8'h0, 8'h59, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h6f, 8'h91, 8'h70, 8'h71, 8'h64, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h2, 8'h3, 8'h2, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h40, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h3e, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h87, 8'h0, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7e, 8'h53, 8'h79, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h54, 8'h0, 8'h0, 8'h0, 8'h23, 8'h53, 8'h62, 8'h10, 8'h0, 8'h27, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h80, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h14, 8'h65, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h5d, 8'h4, 8'h0, 8'h0, 8'h34, 8'h7f, 8'h9b, 8'h9b, 8'h94, 8'h70, 8'h5f, 8'h7b, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h59, 8'h4b, 8'h0, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3f, 8'h0, 8'h3e, 8'h65, 8'h0, 8'h0, 8'h7a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h70, 8'h0, 8'h0, 8'h2, 8'h2, 8'h2, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h71, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h2, 8'h0, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h22, 8'h0, 8'h0, 8'h0, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h3f, 8'h0, 8'h40, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h0, 8'h0, 8'h64, 8'h70, 8'h6f, 8'h70, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h0, 8'h0, 8'h12, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h77, 8'h63, 8'h78, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h51, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h79, 8'h8b, 8'h77, 8'h0, 8'h0, 8'h39, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h81, 8'h50, 8'h28, 8'h37, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h86, 8'h5b, 8'h14, 8'h0, 8'h0, 8'h19, 8'h6c, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h67, 8'h19, 8'h0, 8'h0, 8'h2b, 8'h75, 8'h97, 8'h9b, 8'h92, 8'h72, 8'h5f, 8'h70, 8'h94, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h22, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h2, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h13, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h65, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h23, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h31, 8'h3f, 8'h3f, 8'h3f, 8'h64, 8'h70, 8'h70, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h6f, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h7b, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h0, 8'h0, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h31, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h7a, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h70, 8'h65, 8'h79, 8'h9a, 8'h94, 8'h6d, 8'h17, 8'h0, 8'h0, 8'h35, 8'h7b, 8'h98, 8'h9a, 8'h7a, 8'h0, 8'h0, 8'h2a, 8'h74, 8'h51, 8'h42, 8'h33, 8'h19, 8'h0, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h70, 8'he, 8'h0, 8'h0, 8'h20, 8'h75, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6f, 8'h21, 8'h0, 8'h0, 8'h10, 8'h73, 8'h97, 8'h9a, 8'h94, 8'h7c, 8'h58, 8'h67, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h22, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h3, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h13, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3e, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h85, 8'h9b, 8'h9a, 8'h3f, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h4d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h0, 8'h13, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h31, 8'h0, 8'h3f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h0, 8'h0, 8'h70, 8'h70, 8'h71, 8'h70, 8'h70, 8'h70, 8'h2, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h59, 8'h0, 8'h0, 8'h71, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h66, 8'h5b, 8'h83, 8'h87, 8'h40, 8'h0, 8'h0, 8'h18, 8'h76, 8'h98, 8'h9b, 8'h9b, 8'h82, 8'h1b, 8'h0, 8'h0, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h67, 8'ha, 8'h0, 8'h0, 8'h33, 8'h75, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h76, 8'h25, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h8c, 8'h9a, 8'h97, 8'h84, 8'h59, 8'h5c, 8'h7d, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9a, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h22, 8'h9a, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h2, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h12, 8'h0, 8'h13, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h40, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h13, 8'h9a, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h40, 8'h0, 8'h0, 8'h7c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h58, 8'h0, 8'h0, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h0, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h3e, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7c, 8'h5d, 8'h56, 8'h73, 8'h2d, 8'h0, 8'ha, 8'h79, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h51, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h11, 8'h0, 8'h0, 8'h20, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h5e, 8'h6, 8'h0, 8'h0, 8'h2d, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6d, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h70, 8'h95, 8'h8e, 8'h6c, 8'h4d, 8'h7c, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h2, 8'h0, 8'h71, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h3e, 8'h40, 8'h3f, 8'h3f, 8'h86, 8'h9b, 8'h9b, 8'h91, 8'h4b, 8'h14, 8'h0, 8'h0, 8'h2, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h22, 8'h0, 8'h0, 8'h0, 8'h59, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9a, 8'h87, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h3f, 8'h3d, 8'h40, 8'h31, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h0, 8'h0, 8'h2, 8'h3e, 8'h31, 8'h2, 8'h32, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h6f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h0, 8'h32, 8'h70, 8'h70, 8'h58, 8'h3, 8'h0, 8'h0, 8'h59, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h71, 8'h31, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h2, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h14, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h13, 8'h0, 8'h0, 8'h7b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h1, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h75, 8'h4b, 8'h66, 8'h75, 8'h78, 8'h7f, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h80, 8'h74, 8'h73, 8'h79, 8'h79, 8'h63, 8'h17, 8'h0, 8'h0, 8'h55, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h56, 8'h0, 8'h0, 8'h0, 8'hc, 8'h52, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h6e, 8'h76, 8'h58, 8'h79, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h0, 8'h22, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h21, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h4b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h65, 8'h9a, 8'h9b, 8'h85, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h0, 8'h0, 8'h4c, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h0, 8'h22, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h2, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h4c, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h0, 8'h0, 8'h86, 8'h9b, 8'h9b, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h0, 8'h0, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h72, 8'h56, 8'h75, 8'h93, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h98, 8'h9a, 8'h8a, 8'h3d, 8'h0, 8'h0, 8'h25, 8'h79, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h85, 8'h57, 8'h7, 8'h0, 8'h0, 8'h0, 8'h41, 8'h7f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h7f, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h0, 8'h6, 8'h45, 8'h66, 8'h70, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h64, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h86, 8'h70, 8'h70, 8'h70, 8'h70, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h86, 8'h64, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h86, 8'h64, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6f, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h70, 8'h58, 8'h3f, 8'h4c, 8'h70, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h86, 8'h70, 8'h70, 8'h70, 8'h70, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6f, 8'h6f, 8'h70, 8'h70, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h64, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h86, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h6c, 8'h65, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'h1c, 8'h0, 8'h0, 8'h5f, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8c, 8'h62, 8'h12, 8'h0, 8'h0, 8'h0, 8'h38, 8'h74, 8'h92, 8'h9b, 8'h9a, 8'h89, 8'h49, 8'h0, 8'h0, 8'h10, 8'h44, 8'h0, 8'h0, 8'h18, 8'h0, 8'hd, 8'h3d, 8'h6a, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h69, 8'h66, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h72, 8'h7, 8'h0, 8'h0, 8'h7c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h7a, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h6c, 8'h88, 8'h87, 8'h62, 8'h0, 8'h0, 8'h14, 8'h82, 8'h72, 8'h9, 8'h0, 8'h0, 8'h0, 8'h22, 8'h59, 8'h80, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h85, 8'h63, 8'h5c, 8'h90, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h51, 8'h0, 8'h0, 8'ha, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h81, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h1d, 8'h0, 8'h0, 8'h15, 8'h77, 8'h9a, 8'h8a, 8'h4c, 8'h1, 8'h0, 8'h21, 8'h4f, 8'h7a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h79, 8'h59, 8'h62, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h23, 8'h0, 8'h0, 8'h4c, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h59, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h60, 8'h95, 8'h9a, 8'h97, 8'h81, 8'h62, 8'h46, 8'h4a, 8'h76, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h6f, 8'h50, 8'h77, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h81, 8'h11, 8'h0, 8'h0, 8'h0, 8'hb, 8'h15, 8'h41, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8c, 8'h63, 8'h28, 8'h0, 8'h0, 8'h0, 8'h0, 8'h50, 8'h8a, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h83, 8'h6b, 8'h72, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h89, 8'h67, 8'h60, 8'h81, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h89, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h82, 8'h54, 8'h17, 8'h2, 8'h48, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h72, 8'h6f, 8'h94, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h88, 8'h61, 8'h6d, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6a, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h92, 8'h8b, 8'h88, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h70, 8'h6d, 8'h88, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h60, 8'h67, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h71, 8'h33, 8'h0, 8'h0, 8'h0, 8'h7, 8'h5f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7c, 8'h6b, 8'h77, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h73, 8'h5c, 8'h6a, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h7c, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h64, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h6a, 8'h75, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h66, 8'h52, 8'h81, 8'h94, 8'h9b, 8'h9b, 8'h89, 8'h56, 8'h12, 8'h0, 8'h0, 8'h0, 8'h27, 8'h6a, 8'h8f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8e, 8'h75, 8'h73, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7f, 8'h5f, 8'h62, 8'h8b, 8'h96, 8'h7d, 8'h46, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h78, 8'h92, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h78, 8'h63, 8'h8c, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7e, 8'h59, 8'h77, 8'h88, 8'h52, 8'h0, 8'h0, 8'h0, 8'h11, 8'h58, 8'h8d, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h7b, 8'h66, 8'h7c, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7e, 8'h57, 8'h66, 8'h3b, 8'h0, 8'h0, 8'h30, 8'h74, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h8a, 8'h6d, 8'h6a, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8e, 8'h65, 8'h5a, 8'h5b, 8'h58, 8'h5f, 8'h7f, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h93, 8'h75, 8'h71, 8'h86, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h5e, 8'h60, 8'h88, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h89, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7d, 8'h71, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h75, 8'h61, 8'h73, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h84, 8'h62, 8'h4a, 8'h63, 8'h7a, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h85, 8'h65, 8'h7b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h71, 8'h55, 8'h86, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h43, 8'h0, 8'h0, 8'h0, 8'h10, 8'h61, 8'h94, 8'h97, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h88, 8'h68, 8'h68, 8'h88, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h67, 8'h58, 8'h85, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h33, 8'h79, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7d, 8'h5d, 8'h83, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h7b, 8'h4f, 8'h71, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h69, 8'h39, 8'h49, 8'h71, 8'h92, 8'h99, 8'h8d, 8'h40, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h57, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h82, 8'h72, 8'h7c, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h92, 8'h8d, 8'h8b, 8'h8b, 8'h8e, 8'h94, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h70, 8'h5f, 8'h7b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h7b, 8'h2d, 8'h0, 8'h0, 8'h1a, 8'h3c, 8'h4c, 8'h57, 8'h54, 8'h13, 8'h0, 8'h0, 8'h7, 8'h5, 8'h0, 8'h0, 8'h0, 8'h1, 8'h3a, 8'h6e, 8'h97, 8'h97, 8'h87, 8'h71, 8'h72, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8b, 8'h6b, 8'h30, 8'h0, 8'h0, 8'h0, 8'h12, 8'h8a, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h68, 8'h6a, 8'h88, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h13, 8'h0, 8'h0, 8'h4f, 8'h74, 8'h4e, 8'h4, 8'h0, 8'h0, 8'h0, 8'h14, 8'h71, 8'h87, 8'h71, 8'h6f, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h81, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h80, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h83, 8'h63, 8'h65, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h6b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h80, 8'h90, 8'h75, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h60, 8'h77, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h7a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h89, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h69, 8'h57, 8'h7a, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h51, 8'h0, 8'h0, 8'h0, 8'h41, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h8d, 8'h9b, 8'h94, 8'h79, 8'h43, 8'h0, 8'h0, 8'h0, 8'h3, 8'h5d, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h88, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h8c, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h88, 8'h67, 8'h56, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h84, 8'h31, 8'h0, 8'h0, 8'h71, 8'h65, 8'h3f, 8'h25, 8'h26, 8'h36, 8'h77, 8'h97, 8'h9a, 8'h9b, 8'h97, 8'h84, 8'h51, 8'hd, 8'h0, 8'h17, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h72, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h78, 8'h9a, 8'h99, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h80, 8'h60, 8'h6e, 8'h8d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h64, 8'he, 8'h0, 8'h5b, 8'h88, 8'h90, 8'h8e, 8'h8b, 8'h8d, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8b, 8'h5d, 8'h27, 8'h5c, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h83, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h93, 8'h87, 8'h7d, 8'h89, 8'h96, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h79, 8'h54, 8'h78, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8f, 8'h86, 8'h86, 8'h84, 8'h6e, 8'h19, 8'h0, 8'h38, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h71, 8'h62, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h13, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h81, 8'h5c, 8'h0, 8'h53, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h5b, 8'h64, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h55, 8'h21, 8'h21, 8'h1b, 8'hd, 8'h0, 8'h0, 8'h31, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h6a, 8'h5f, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'he, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h75, 8'h1b, 8'h0, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h83, 8'h58, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h63, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h74, 8'h5e, 8'h71, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7d, 8'h30, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h78, 8'h1f, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h93, 8'h72, 8'h62, 8'h75, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h18, 8'h0, 8'h0, 8'ha, 8'h14, 8'h13, 8'h1d, 8'h43, 8'h87, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h5f, 8'h66, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h7e, 8'h40, 8'h0, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h63, 8'h5e, 8'h91, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h29, 8'h0, 8'h0, 8'h26, 8'h33, 8'h36, 8'h40, 8'h63, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h76, 8'h63, 8'h7a, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h72, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h75, 8'h83, 8'h49, 8'h0, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h75, 8'h5e, 8'h71, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h6d, 8'h16, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h72, 8'h8c, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h7e, 8'h53, 8'h7a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h5e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h55, 8'h90, 8'h86, 8'h56, 8'h0, 8'h0, 8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h70, 8'h4c, 8'h85, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h70, 8'h29, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h7d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h83, 8'h5f, 8'h58, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h8f, 8'h9a, 8'h8b, 8'h63, 8'h0, 8'h0, 8'h0, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h83, 8'h5c, 8'h5f, 8'h86, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h78, 8'h4c, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h45, 8'h84, 8'h99, 8'h9b, 8'h95, 8'h74, 8'h50, 8'h7c, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h81, 8'h63, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h66, 8'h7f, 8'h8b, 8'h85, 8'h75, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h97, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h78, 8'h52, 8'h7b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h90, 8'h67, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h49, 8'h7a, 8'h7b, 8'h64, 8'h68, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h83, 8'h47, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h7f, 8'h77, 8'h5d, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8e, 8'h6a, 8'h6a, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7d, 8'h8, 8'h0, 8'h15, 8'h59, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h43, 8'h50, 8'h8a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h69, 8'h0, 8'h0, 8'h3, 8'h46, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h5d, 8'h69, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h95, 8'h91, 8'h95, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7f, 8'ha, 8'h0, 8'ha, 8'h8b, 8'h80, 8'h50, 8'hb, 8'h0, 8'h0, 8'h0, 8'h8, 8'h43, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8c, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h40, 8'h6a, 8'h67, 8'h73, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h69, 8'h5e, 8'h7a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8a, 8'h63, 8'h3f, 8'h5f, 8'h87, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7f, 8'h9, 8'h0, 8'h0, 8'h8e, 8'h99, 8'h8d, 8'h7a, 8'h69, 8'h52, 8'h36, 8'h55, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h8b, 8'h79, 8'h57, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h33, 8'h54, 8'h66, 8'h7e, 8'h93, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h63, 8'h5c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h59, 8'h0, 8'h0, 8'h0, 8'h8, 8'h1f, 8'h44, 8'h7c, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h18, 8'h0, 8'h0, 8'h8a, 8'h9b, 8'h9a, 8'h98, 8'h8b, 8'h68, 8'h58, 8'h79, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h8e, 8'h7c, 8'h5b, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4a, 8'h83, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h78, 8'h60, 8'h6f, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h35, 8'h3c, 8'h40, 8'h44, 8'h34, 8'h0, 8'h0, 8'h0, 8'h78, 8'h95, 8'h9b, 8'h99, 8'h84, 8'h56, 8'h6e, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h8b, 8'h74, 8'h29, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h64, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h6b, 8'h51, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7d, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h91, 8'h99, 8'h8e, 8'h72, 8'h54, 8'h82, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'h33, 8'h0, 8'h0, 8'h0, 8'h0, 8'ha, 8'h2, 8'h0, 8'h0, 8'h84, 8'h96, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7b, 8'h55, 8'h7b, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h85, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5, 8'h87, 8'h98, 8'h95, 8'h74, 8'h54, 8'h78, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h9, 8'h56, 8'h69, 8'h2, 8'h0, 8'h0, 8'h91, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7f, 8'h56, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h50, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h63, 8'h61, 8'h5b, 8'h58, 8'h59, 8'h59, 8'h5e, 8'h74, 8'h97, 8'h9a, 8'h91, 8'h6b, 8'h51, 8'h8e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h80, 8'h7, 8'h0, 8'h0, 8'h54, 8'h85, 8'h92, 8'h7d, 8'h0, 8'h0, 8'h0, 8'h97, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8a, 8'h58, 8'h6d, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h98, 8'h83, 8'h45, 8'h0, 8'h0, 8'h14, 8'h6b, 8'h96, 8'h94, 8'h90, 8'h92, 8'h92, 8'h93, 8'h96, 8'h9a, 8'h95, 8'h76, 8'h66, 8'h7a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h67, 8'h0, 8'h0, 8'h23, 8'h85, 8'h99, 8'h91, 8'h72, 8'h0, 8'h0, 8'h0, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h77, 8'h62, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7d, 8'h38, 8'h0, 8'h0, 8'h2a, 8'h78, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h61, 8'h66, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8a, 8'h52, 8'h0, 8'h0, 8'h41, 8'h8b, 8'h9b, 8'h8c, 8'h6b, 8'h0, 8'h0, 8'h1, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8d, 8'h63, 8'h62, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h73, 8'h20, 8'h0, 8'h0, 8'h44, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h74, 8'h62, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h84, 8'h41, 8'h0, 8'h0, 8'h64, 8'h92, 8'h9b, 8'h89, 8'h5d, 8'h0, 8'h0, 8'h15, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h75, 8'h5e, 8'h6a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h6a, 8'h0, 8'h0, 8'h25, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h56, 8'h70, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7b, 8'h20, 8'h0, 8'h0, 8'h8b, 8'h98, 8'h9a, 8'h84, 8'h4a, 8'h0, 8'h0, 8'h36, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h68, 8'h57, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h34, 8'h0, 8'h0, 8'h52, 8'h99, 8'h9b, 8'h9b, 8'h99, 8'h8d, 8'h69, 8'h5a, 8'h7d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h66, 8'h0, 8'h0, 8'h0, 8'h97, 8'h9a, 8'h9b, 8'h7e, 8'h37, 8'h0, 8'h0, 8'h38, 8'h96, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h80, 8'h62, 8'h64, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h4c, 8'h0, 8'h0, 8'h3f, 8'h98, 8'h9b, 8'h9b, 8'h99, 8'h7e, 8'h51, 8'h71, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h5b, 8'h0, 8'h0, 8'h21, 8'h9a, 8'h9b, 8'h9b, 8'h7e, 8'h35, 8'h0, 8'h0, 8'h43, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h6f, 8'h4e, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h7a, 8'h1e, 8'h0, 8'h0, 8'h5e, 8'h99, 8'h9b, 8'h99, 8'h8b, 8'h6c, 8'h54, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h61, 8'h0, 8'h0, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h2e, 8'h0, 8'h0, 8'h56, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h84, 8'h5e, 8'h73, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h89, 8'h6f, 8'h3c, 8'h0, 8'h0, 8'h30, 8'h8e, 8'h9a, 8'h9b, 8'h96, 8'h75, 8'h5a, 8'h74, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8f, 8'h7b, 8'h51, 8'h34, 8'h87, 8'h9b, 8'h9b, 8'h9a, 8'h7d, 8'h1f, 8'h0, 8'h0, 8'h6c, 8'h98, 8'h98, 8'h98, 8'h96, 8'h97, 8'h93, 8'h93, 8'h93, 8'h93, 8'h95, 8'h98, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7f, 8'h5a, 8'h78, 8'h99, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h48, 8'h0, 8'h0, 8'h0, 8'h25, 8'h78, 8'h9a, 8'h9b, 8'h9b, 8'h93, 8'h6b, 8'h51, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h94, 8'h8e, 8'h92, 8'h97, 8'h9b, 8'h9b, 8'h97, 8'h79, 8'h0, 8'h0, 8'h0, 8'h65, 8'h75, 8'h76, 8'h75, 8'h72, 8'h6e, 8'h6a, 8'h68, 8'h67, 8'h69, 8'h6f, 8'h79, 8'h88, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8b, 8'h56, 8'h6f, 8'h91, 8'h9a, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h75, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h6b, 8'h93, 8'h9b, 8'h9a, 8'h93, 8'h74, 8'h63, 8'h77, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h0, 8'h7, 8'h22, 8'h3d, 8'h82, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7c, 8'h63, 8'h73, 8'h9b, 8'h9a, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7e, 8'h4f, 8'hb, 8'h0, 8'h0, 8'h0, 8'ha, 8'h38, 8'h6d, 8'h8f, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h63, 8'h63, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h81, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h61, 8'h63, 8'h91, 8'h99, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h69, 8'h8f, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h7a, 8'h64, 8'h75, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h60, 8'h54, 8'h57, 8'h58, 8'h42, 8'h34, 8'h2f, 8'h37, 8'h2e, 8'h53, 8'h8, 8'h0, 8'h0, 8'h0, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h73, 8'h62, 8'h75, 8'h99, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h2e, 8'h0, 8'h0, 8'h0, 8'h31, 8'h6e, 8'h88, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8b, 8'h58, 8'h6f, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h92, 8'h73, 8'hb, 8'h0, 8'h0, 8'h29, 8'h73, 8'h8b, 8'h87, 8'h88, 8'h8a, 8'h8b, 8'h8e, 8'h91, 8'h94, 8'h97, 8'h99, 8'h69, 8'ha, 8'h0, 8'h0, 8'h76, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h99, 8'h99, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h99, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h69, 8'h55, 8'h91, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h72, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h84, 8'h53, 8'h76, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h7d, 8'h32, 8'h0, 8'h0, 8'h1a, 8'h75, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h11, 8'h0, 8'h0, 8'h65, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h94, 8'h92, 8'h91, 8'h90, 8'h90, 8'h8c, 8'h87, 8'h83, 8'h7b, 8'h71, 8'h68, 8'h60, 8'h5f, 8'h5f, 8'h5d, 8'h5c, 8'h5d, 8'h5f, 8'h5f, 8'h63, 8'h65, 8'h6a, 8'h72, 8'h78, 8'h7d, 8'h84, 8'h8b, 8'h8e, 8'h90, 8'h91, 8'h93, 8'h94, 8'h96, 8'h98, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h74, 8'h56, 8'h80, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h76, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h44, 8'h7d, 8'h95, 8'h82, 8'h5d, 8'h73, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h83, 8'h55, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h33, 8'h0, 8'h0, 8'h4a, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h95, 8'h92, 8'h90, 8'h8e, 8'h87, 8'h78, 8'h5d, 8'h37, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h35, 8'h53, 8'h6c, 8'h7f, 8'h8b, 8'h90, 8'h92, 8'h95, 8'h96, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8a, 8'h6e, 8'h59, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h86, 8'h54, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h5e, 8'h69, 8'h4a, 8'h85, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h60, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h61, 8'h0, 8'h0, 8'h20, 8'h94, 8'h9a, 8'h9b, 8'h98, 8'h95, 8'h90, 8'h82, 8'h5b, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h41, 8'h6f, 8'h87, 8'h90, 8'h92, 8'h95, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h7d, 8'h4f, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h93, 8'h80, 8'h47, 8'h5, 8'h0, 8'h0, 8'h0, 8'h24, 8'h3b, 8'h52, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h92, 8'h61, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h76, 8'h0, 8'h0, 8'h0, 8'h6e, 8'h7c, 8'h85, 8'h69, 8'h13, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h2f, 8'h4d, 8'h62, 8'h72, 8'h7e, 8'h89, 8'h8f, 8'h94, 8'h97, 8'h96, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h93, 8'h8e, 8'h87, 8'h81, 8'h76, 8'h66, 8'h51, 8'h3d, 8'h25, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h5e, 8'h80, 8'h8f, 8'h92, 8'h97, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8a, 8'h64, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h8f, 8'h7c, 8'h54, 8'h29, 8'h3a, 8'h1c, 8'h6, 8'h65, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h6d, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h7e, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h82, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h9, 8'h1a, 8'h2d, 8'h48, 8'h69, 8'h84, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h88, 8'h6e, 8'h49, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h64, 8'h86, 8'h91, 8'h93, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h86, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h90, 8'h86, 8'h7d, 8'h55, 8'h46, 8'h8f, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h80, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h97, 8'h95, 8'h95, 8'h93, 8'h91, 8'h91, 8'h91, 8'h90, 8'h8f, 8'h90, 8'h91, 8'h91, 8'h90, 8'h91, 8'h92, 8'h93, 8'h94, 8'h96, 8'h96, 8'h98, 8'h9a, 8'h98, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h89, 8'h67, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h5b, 8'h86, 8'h91, 8'h95, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h6c, 8'h66, 8'h81, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h2f, 8'h0, 8'h0, 8'h11, 8'h72, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h38, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h92, 8'h91, 8'h8f, 8'h90, 8'h8f, 8'h8e, 8'h8c, 8'h82, 8'h6d, 8'h53, 8'h37, 8'h1d, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h29, 8'h49, 8'h60, 8'h69, 8'h4f, 8'h65, 8'h8f, 8'h8f, 8'h8f, 8'h90, 8'h93, 8'h94, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h70, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h6b, 8'h89, 8'h95, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h5f, 8'h69, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8b, 8'h35, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h8f, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h8e, 8'h6f, 8'h5a, 8'h53, 8'h66, 8'h81, 8'h92, 8'h98, 8'h93, 8'h90, 8'h8f, 8'h8f, 8'h8a, 8'h73, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6, 8'h3, 8'h2, 8'h5, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h13, 8'h53, 8'h81, 8'h8f, 8'h8f, 8'h90, 8'h90, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h82, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4f, 8'h85, 8'h92, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h7a, 8'h65, 8'h78, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h6b, 8'h0, 8'h0, 8'h0, 8'h47, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h96, 8'h8f, 8'h8f, 8'h8f, 8'h83, 8'h4f, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h35, 8'h6c, 8'h8a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h59, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4, 8'h69, 8'h93, 8'h7c, 8'h52, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h6b, 8'h8a, 8'h90, 8'h90, 8'h93, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7f, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h7f, 8'h91, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h58, 8'h75, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h8b, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h7f, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h90, 8'h8e, 8'h7c, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h5b, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h8e, 8'h26, 8'h0, 8'h0, 8'h0, 8'hb, 8'h56, 8'h86, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h7b, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h88, 8'h8e, 8'h91, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h71, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h7e, 8'h94, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h52, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h7c, 8'h0, 8'h0, 8'h0, 8'h74, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h93, 8'h8f, 8'h8c, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h47, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h77, 8'h7, 8'h0, 8'h0, 8'h24, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h65, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h77, 8'h8f, 8'h90, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h84, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h87, 8'h94, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h82, 8'h60, 8'h6e, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h7f, 8'h0, 8'h0, 8'h0, 8'h71, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h91, 8'h8d, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h41, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h7c, 8'h8e, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h64, 8'h8d, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h75, 8'h49, 8'h84, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h90, 8'h74, 8'h31, 8'h1b, 8'h0, 8'h0, 8'h54, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h95, 8'h8e, 8'h7a, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h86, 8'h1c, 8'h0, 8'h0, 8'h1, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h5e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4f, 8'h8c, 8'h90, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7f, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h80, 8'h95, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h6d, 8'h54, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h7e, 8'h21, 8'h0, 8'h0, 8'h0, 8'h20, 8'h0, 8'h0, 8'h3a, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h8f, 8'h6a, 8'h5, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h7a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h64, 8'h0, 8'h0, 8'h0, 8'h34, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8e, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h84, 8'h90, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6c, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'ha, 8'h6a, 8'h90, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h72, 8'h5c, 8'h7b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h90, 8'h63, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h85, 8'h8d, 8'h4e, 8'h36, 8'h73, 8'h8e, 8'h99, 8'h93, 8'h8f, 8'h6a, 8'h2, 8'h0, 8'h0, 8'h0, 8'h3f, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h93, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h67, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h6, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h82, 8'h90, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h8a, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h68, 8'h59, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8e, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h8e, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h95, 8'h8f, 8'h8e, 8'h6c, 8'h5, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h70, 8'h2, 8'h0, 8'h0, 8'h13, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7e, 8'h14, 8'h0, 8'h0, 8'h0, 8'h33, 8'h88, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h73, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h82, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7c, 8'h62, 8'h6b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h84, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h91, 8'h85, 8'h2d, 8'h0, 8'h0, 8'h0, 8'h48, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8d, 8'h35, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h8f, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h87, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h79, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h66, 8'h63, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h7f, 8'h22, 8'h0, 8'h0, 8'h0, 8'h0, 8'h69, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h90, 8'h5a, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h87, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h52, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h7d, 8'h92, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8c, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h78, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h87, 8'h5a, 8'h6b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7a, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h68, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h88, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8e, 8'h28, 8'h0, 8'h0, 8'h0, 8'h55, 8'h90, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h46, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h79, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h73, 8'h5e, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h99, 8'h96, 8'h80, 8'h20, 8'h0, 8'h0, 8'h0, 8'h2, 8'h6d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h91, 8'h77, 8'hb, 8'h0, 8'h0, 8'h29, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h78, 8'h6, 8'h0, 8'h0, 8'h2f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h61, 8'h0, 8'h0, 8'h0, 8'h36, 8'h8e, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h7b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h59, 8'h74, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h86, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h92, 8'h5a, 8'h0, 8'h0, 8'h0, 8'h4f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h78, 8'h15, 8'h0, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h19, 8'h0, 8'h0, 8'h19, 8'h7f, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h87, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h80, 8'h52, 8'h7d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h62, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h91, 8'h46, 8'h0, 8'h0, 8'h1, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h73, 8'ha, 8'h0, 8'h0, 8'h0, 8'h22, 8'h88, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h34, 8'h0, 8'h0, 8'hb, 8'h75, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h48, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h90, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h89, 8'h6b, 8'h67, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h94, 8'h64, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h91, 8'h41, 8'h0, 8'h0, 8'h15, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h95, 8'h91, 8'h8f, 8'h8e, 8'h90, 8'h8f, 8'h91, 8'h94, 8'h99, 8'h94, 8'h7f, 8'h15, 8'h0, 8'h0, 8'h0, 8'h30, 8'h8c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h43, 8'h0, 8'h0, 8'h5, 8'h72, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h42, 8'h0, 8'h0, 8'h0, 8'h0, 8'h61, 8'h94, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h76, 8'h50, 8'h86, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7b, 8'h15, 8'h0, 8'h0, 8'h0, 8'h39, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h41, 8'h0, 8'h0, 8'h1c, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h85, 8'h66, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h57, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h29, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h0, 8'h6, 8'h73, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h13, 8'h7a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h71, 8'h4a, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h8f, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h91, 8'h49, 8'h0, 8'h0, 8'h1d, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h93, 8'h7b, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h0, 8'hf, 8'h79, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h79, 8'hd, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h90, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h7c, 8'h67, 8'h6f, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h66, 8'h0, 8'h0, 8'h0, 8'h6, 8'h73, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h5e, 8'h0, 8'h0, 8'h12, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h67, 8'h94, 8'h97, 8'h97, 8'h8e, 8'h63, 8'h19, 8'h0, 8'h11, 8'h69, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h46, 8'h0, 8'h0, 8'h1e, 8'h86, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h63, 8'h95, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h6b, 8'h5e, 8'h8d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h8e, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h50, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h75, 8'h9, 8'h0, 8'hc, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h94, 8'h61, 8'h0, 8'h0, 8'h0, 8'h0, 8'h9, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h39, 8'h0, 8'h0, 8'h30, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h38, 8'h0, 8'h0, 8'h0, 8'h25, 8'h88, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h88, 8'h62, 8'h60, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h61, 8'h0, 8'h0, 8'h0, 8'h28, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h8a, 8'h22, 8'h0, 8'h0, 8'h5e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h93, 8'h61, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h27, 8'h0, 8'h0, 8'h53, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h13, 8'h0, 8'h0, 8'h0, 8'h5f, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h74, 8'h63, 8'h72, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h23, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h37, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h78, 8'h11, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h80, 8'h11, 8'h0, 8'hc, 8'h78, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h53, 8'h0, 8'h0, 8'h0, 8'h24, 8'h87, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8d, 8'h5e, 8'h6d, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h6b, 8'h0, 8'h0, 8'h0, 8'h35, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h68, 8'h0, 8'h0, 8'h28, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h71, 8'h8, 8'h0, 8'h0, 8'h0, 8'h29, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h56, 8'h0, 8'h0, 8'h2b, 8'h91, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h62, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h5a, 8'h6e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h93, 8'h32, 8'h0, 8'h0, 8'h7, 8'h77, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h8f, 8'h24, 8'h0, 8'h0, 8'h6a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h94, 8'h38, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h0, 8'h52, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h92, 8'h72, 8'h69, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h84, 8'h12, 8'h0, 8'h0, 8'h36, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h4e, 8'h0, 8'h0, 8'h3c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h81, 8'h13, 8'h0, 8'h0, 8'h1c, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hf, 8'h0, 8'h1c, 8'h88, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h1c, 8'h0, 8'h0, 8'h8, 8'h77, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h56, 8'h7a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h62, 8'h0, 8'h0, 8'h0, 8'h6a, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h8b, 8'h1c, 8'h0, 8'h13, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h46, 8'h0, 8'h0, 8'h44, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h51, 8'h0, 8'h0, 8'h0, 8'h48, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h7d, 8'h4e, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h40, 8'h0, 8'h0, 8'h3b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h51, 8'h0, 8'h0, 8'h44, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h94, 8'h8f, 8'h91, 8'h97, 8'h9b, 8'h95, 8'h3b, 8'h0, 8'h0, 8'h15, 8'h82, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h1d, 8'h0, 8'h1b, 8'h89, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h12, 8'h0, 8'h0, 8'h26, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8a, 8'h6b, 8'h5c, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h93, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8f, 8'h28, 8'h0, 8'h0, 8'h67, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h23, 8'h0, 8'h12, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h58, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h8c, 8'h31, 8'h0, 8'h0, 8'h31, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h49, 8'h0, 8'h0, 8'h4d, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h36, 8'h0, 8'h0, 8'hc, 8'h7e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h77, 8'h57, 8'h7e, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h91, 8'h8c, 8'h91, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7f, 8'h15, 8'h0, 8'h29, 8'h8c, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h69, 8'h0, 8'h0, 8'h3b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h7d, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h33, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h86, 8'h15, 8'h0, 8'h28, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h63, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6f, 8'h4d, 8'h8e, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h63, 8'h0, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h30, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h92, 8'h91, 8'h8b, 8'h68, 8'h2c, 8'h0, 8'h0, 8'h0, 8'h42, 8'h98, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h4b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3b, 8'h0, 8'h0, 8'h6c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h20, 8'h0, 8'h0, 8'h5c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8c, 8'h6a, 8'h58, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h48, 8'h0, 8'h6, 8'h6f, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h88, 8'h17, 8'h0, 8'h2d, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h91, 8'h92, 8'h91, 8'h90, 8'h88, 8'h4c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h8d, 8'h9a, 8'h9b, 8'h92, 8'h50, 8'h49, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h66, 8'h0, 8'h0, 8'h36, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h54, 8'h0, 8'h0, 8'h47, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h75, 8'h64, 8'h7c, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h39, 8'h0, 8'h2a, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h59, 8'h0, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h59, 8'h8a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h1f, 8'h0, 8'h1d, 8'h8d, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h79, 8'hf, 8'h0, 8'h3c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h64, 8'h5f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h2d, 8'h0, 8'h43, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h31, 8'h0, 8'hd, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h3c, 8'h0, 8'h0, 8'h8, 8'h4, 8'h2e, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h39, 8'h0, 8'h0, 8'h71, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h33, 8'h0, 8'h3a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h63, 8'h63, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h21, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h1e, 8'h0, 8'h2d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3d, 8'h0, 8'h0, 8'h2b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5f, 8'h0, 8'h0, 8'h40, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h3a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h78, 8'h6b, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7c, 8'h1a, 8'h11, 8'h72, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h7d, 8'hc, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h19, 8'h0, 8'h2a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h17, 8'h0, 8'h29, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h72, 8'h1f, 8'h42, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h60, 8'h70, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h70, 8'h12, 8'h24, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h54, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h42, 8'h0, 8'h0, 8'h63, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h2c, 8'h0, 8'h1b, 8'h8d, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h89, 8'h48, 8'h56, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h56, 8'h6f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h5e, 8'h8, 8'h37, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h39, 8'h0, 8'h14, 8'h85, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h79, 8'h4, 8'h0, 8'h2e, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h98, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3a, 8'h0, 8'h8, 8'h7a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h98, 8'h85, 8'h59, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h59, 8'h6, 8'h45, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h28, 8'h0, 8'h27, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h96, 8'h93, 8'h5d, 8'h0, 8'h0, 8'hb, 8'h7c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h81, 8'h67, 8'h5d, 8'h68, 8'h81, 8'h8f, 8'h92, 8'h97, 8'h95, 8'h91, 8'h90, 8'h8f, 8'h8f, 8'h8f, 8'h8f, 8'h8f, 8'h91, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h56, 8'h0, 8'h0, 8'h5b, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h8b, 8'h67, 8'h70, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h5d, 8'h15, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h20, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h96, 8'h92, 8'h8b, 8'h64, 8'h34, 8'h0, 8'h0, 8'h0, 8'h9, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h95, 8'h96, 8'h98, 8'h97, 8'h97, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h84, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h33, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h48, 8'h8d, 8'h99, 8'h9b, 8'h9a, 8'h97, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h74, 8'h0, 8'h0, 8'h40, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h99, 8'h82, 8'h50, 8'h7e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h53, 8'hd, 8'h51, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h8f, 8'h18, 8'h0, 8'h3c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h91, 8'h72, 8'h34, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h89, 8'h99, 8'h94, 8'h89, 8'h8c, 8'h9a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h90, 8'h5f, 8'h36, 8'h3a, 8'h43, 8'h43, 8'h42, 8'h53, 8'h77, 8'h8a, 8'h8d, 8'h78, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h1, 8'h38, 8'h5, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h61, 8'h90, 8'h81, 8'h42, 8'h3b, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h86, 8'h10, 8'h0, 8'h2f, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h97, 8'h7c, 8'h4d, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h4e, 8'hb, 8'h56, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'hf, 8'h0, 8'h47, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h90, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h55, 8'h86, 8'h9a, 8'h94, 8'h69, 8'h17, 8'h0, 8'h20, 8'h6c, 8'h89, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h78, 8'ha, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h7d, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h7f, 8'h5c, 8'h5e, 8'h84, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h28, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h21, 8'h0, 8'h27, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9a, 8'h90, 8'h76, 8'h5b, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h54, 8'h16, 8'h5a, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h79, 8'h5, 8'h0, 8'h56, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h66, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h58, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h1f, 8'h0, 8'h30, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h86, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h49, 8'h4e, 8'h50, 8'h4c, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h25, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h28, 8'h0, 8'h23, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h96, 8'h7a, 8'h5e, 8'h7d, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h5a, 8'h24, 8'h62, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h71, 8'h0, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h75, 8'hf, 8'h0, 8'h0, 8'h0, 8'h46, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h26, 8'h12, 8'h76, 8'h9b, 8'h90, 8'h87, 8'h68, 8'h2, 8'h0, 8'h6e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h56, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h92, 8'h99, 8'h9b, 8'h52, 8'h0, 8'h24, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h2c, 8'h0, 8'h20, 8'h96, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h94, 8'h6e, 8'h52, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h5b, 8'h20, 8'h5e, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h6b, 8'h0, 8'h0, 8'h71, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h69, 8'h2, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h85, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h38, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h65, 8'h96, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h8c, 8'h20, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h15, 8'h0, 8'h74, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h2d, 8'h0, 8'h1d, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h93, 8'h6d, 8'h52, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h73, 8'h48, 8'h6e, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h60, 8'h0, 8'h0, 8'h76, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h82, 8'h18, 8'h0, 8'h0, 8'h0, 8'h10, 8'h79, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h77, 8'ha, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2a, 8'h0, 8'h1a, 8'h36, 8'h59, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h8d, 8'h8a, 8'h8a, 8'h8c, 8'h8f, 8'h93, 8'h96, 8'h96, 8'h97, 8'h99, 8'h98, 8'h92, 8'h8c, 8'h40, 8'h0, 8'h0, 8'h0, 8'h36, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h34, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h8f, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2f, 8'h0, 8'h1c, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h92, 8'h6d, 8'h66, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7e, 8'h5a, 8'h75, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h63, 8'h0, 8'h0, 8'h0, 8'h53, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8b, 8'h44, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h39, 8'h0, 8'h56, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h36, 8'h53, 8'h75, 8'h50, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h54, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h61, 8'h0, 8'h9, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h19, 8'h0, 8'hd, 8'h7d, 8'h96, 8'h98, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h31, 8'h0, 8'h1e, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h8d, 8'h65, 8'h8c, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h85, 8'h63, 8'h78, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h73, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h10, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2c, 8'h0, 8'h52, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h52, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2c, 8'h0, 8'h2d, 8'h91, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h61, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h71, 8'h86, 8'h86, 8'h84, 8'h84, 8'h86, 8'h1d, 8'h0, 8'he, 8'h8a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h8b, 8'h63, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h66, 8'h76, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h6d, 8'h0, 8'h9, 8'h29, 8'h0, 8'h13, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8f, 8'h75, 8'h11, 8'h0, 8'h0, 8'h0, 8'h4f, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h28, 8'h24, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h53, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h2e, 8'h0, 8'h0, 8'h3c, 8'h98, 8'h9a, 8'h99, 8'h8a, 8'h5c, 8'h3d, 8'h3a, 8'h6, 8'h0, 8'h0, 8'h55, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h0, 8'h0, 8'h9, 8'h6b, 8'h95, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h93, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h8c, 8'h8e, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h30, 8'h0, 8'h9, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h8c, 8'h67, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h70, 8'h76, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h77, 8'h2, 8'h3, 8'h76, 8'h23, 8'h0, 8'h29, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8e, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h33, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h28, 8'h21, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h75, 8'h51, 8'h4b, 8'h1b, 8'h0, 8'h31, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h38, 8'h0, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h86, 8'h63, 8'h5f, 8'h82, 8'h92, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h73, 8'hd, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h5d, 8'h89, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h63, 8'hf, 8'h33, 8'h86, 8'h99, 8'h9b, 8'h9a, 8'h95, 8'h88, 8'h1d, 8'h0, 8'h0, 8'h44, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2c, 8'h0, 8'h27, 8'h9b, 8'h7f, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h15, 8'h0, 8'h21, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h91, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h7b, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h8, 8'h0, 8'h6c, 8'h8b, 8'h14, 8'h0, 8'h42, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7f, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h24, 8'h1e, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h7f, 8'h1f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h76, 8'h0, 8'h0, 8'h32, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h10, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h55, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h31, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'hf, 8'h0, 8'h0, 8'h1, 8'h6d, 8'h8f, 8'h81, 8'h27, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h52, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h25, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h97, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h79, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h14, 8'h0, 8'h59, 8'h9a, 8'h84, 8'hc, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h57, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h20, 8'h1a, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h48, 8'h0, 8'h0, 8'h35, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h22, 8'h0, 8'h1a, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h21, 8'h0, 8'h11, 8'h7d, 8'h88, 8'h54, 8'h0, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h8b, 8'h55, 8'h0, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h7a, 8'h2b, 8'h0, 8'h0, 8'h55, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h32, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h29, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h7c, 8'h7a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h19, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h5c, 8'h0, 8'h5, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h88, 8'h2d, 8'h0, 8'h0, 8'h1e, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h21, 8'h1b, 8'h8b, 8'h9b, 8'h99, 8'h8e, 8'h30, 8'h0, 8'h16, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h45, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h5c, 8'h0, 8'h19, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h3d, 8'h0, 8'h24, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h36, 8'h0, 8'h5a, 8'h92, 8'h34, 8'h0, 8'h0, 8'h0, 8'h18, 8'h7d, 8'h9b, 8'h9b, 8'h8e, 8'h1f, 8'h0, 8'h0, 8'h38, 8'h8a, 8'h94, 8'h9a, 8'h9b, 8'h2c, 8'h0, 8'h28, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h25, 8'h0, 8'h32, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h84, 8'h7d, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h1d, 8'h0, 8'h40, 8'h9a, 8'h9a, 8'h9b, 8'h46, 8'h0, 8'h1a, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h50, 8'h0, 8'h0, 8'h0, 8'h35, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h21, 8'h15, 8'h82, 8'h90, 8'h6d, 8'h5, 8'h0, 8'h2c, 8'h8f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h92, 8'h90, 8'h8f, 8'h8c, 8'h89, 8'h89, 8'h39, 8'h0, 8'h0, 8'h2d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h96, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h27, 8'h0, 8'h36, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h46, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h0, 8'h59, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h24, 8'h17, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h93, 8'h27, 8'h0, 8'h0, 8'h0, 8'h20, 8'h7e, 8'h93, 8'h20, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h1c, 8'h0, 8'h42, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h8b, 8'h81, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h24, 8'h0, 8'h37, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h17, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h16, 8'h84, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h24, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h91, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h29, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h8f, 8'h81, 8'h49, 8'h23, 8'h52, 8'h81, 8'h89, 8'h8d, 8'h77, 8'h8, 8'h7, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h14, 8'h0, 8'h3a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h21, 8'h0, 8'h2d, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h78, 8'h4, 8'h2a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h1, 8'h0, 8'h0, 8'h0, 8'h6, 8'h0, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h85, 8'hb, 8'h0, 8'h5a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h81, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h31, 8'h0, 8'h2f, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h1f, 8'h94, 8'h9b, 8'h9a, 8'h8d, 8'h28, 8'h0, 8'h0, 8'h1d, 8'h84, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7a, 8'h52, 8'h49, 8'h48, 8'h66, 8'h8e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8c, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h32, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h9a, 8'h9a, 8'h9b, 8'h96, 8'h20, 8'h0, 8'h23, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6b, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h2f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h89, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h22, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h71, 8'h0, 8'h0, 8'h78, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h47, 8'h0, 8'h29, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h25, 8'h0, 8'h28, 8'h9b, 8'h99, 8'h89, 8'h1b, 8'h0, 8'h5, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h8f, 8'h52, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h6b, 8'h37, 8'h8, 8'h1c, 8'h2, 8'h0, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9a, 8'h37, 8'h0, 8'h0, 8'h67, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h25, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h30, 8'h0, 8'h46, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h5b, 8'h8, 8'h24, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h4e, 8'h0, 8'h15, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h1c, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h28, 8'h95, 8'h67, 8'h0, 8'h0, 8'h3a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h54, 8'h0, 8'h0, 8'h0, 8'h32, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h54, 8'h0, 8'h21, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6c, 8'h0, 8'h0, 8'h2f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h0, 8'h2d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h83, 8'h14, 8'ha, 8'h7d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h38, 8'h0, 8'h1f, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h87, 8'h87, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h11, 8'h0, 8'h77, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h23, 8'h0, 8'h17, 8'h25, 8'h0, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h4e, 8'h0, 8'h0, 8'h2d, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h62, 8'h0, 8'h26, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h79, 8'h0, 8'h0, 8'h19, 8'h8d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h0, 8'h28, 8'h95, 8'h96, 8'h95, 8'h97, 8'h92, 8'h64, 8'he, 8'h0, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h28, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h82, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h1d, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h71, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h43, 8'h0, 8'h28, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h2b, 8'h0, 8'h0, 8'h1d, 8'h2f, 8'h32, 8'h33, 8'h0, 8'h0, 8'h0, 8'h0, 8'h62, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h23, 8'h0, 8'h41, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h89, 8'h8a, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h26, 8'h0, 8'h39, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8b, 8'h14, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h1e, 8'h0, 8'h38, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2d, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'hd, 8'h0, 8'h0, 8'h5e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h14, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h89, 8'hf, 8'h0, 8'h71, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h43, 8'h0, 8'h2c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h42, 8'h2f, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h62, 8'h0, 8'h20, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2f, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'hf, 8'h0, 8'h0, 8'h51, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h7a, 8'h5d, 8'h64, 8'h6b, 8'h79, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h5b, 8'h0, 8'h17, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h75, 8'h0, 8'h20, 8'h92, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h27, 8'h0, 8'h46, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h1b, 8'h0, 8'h35, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h17, 8'h0, 8'h0, 8'h43, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h91, 8'h90, 8'h91, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h1f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h93, 8'h19, 8'h0, 8'h69, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6f, 8'h0, 8'h26, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h33, 8'h0, 8'h0, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h27, 8'h0, 8'h0, 8'h34, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h42, 8'h0, 8'h0, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h27, 8'h0, 8'h33, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h24, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h3b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h4c, 8'h0, 8'h0, 8'h33, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h3c, 8'h0, 8'h0, 8'h1c, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h39, 8'h0, 8'h24, 8'h5e, 8'h1, 8'h2c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h19, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h4a, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'hc, 8'h7, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h92, 8'h90, 8'h8f, 8'h81, 8'h23, 8'h0, 8'h0, 8'h2a, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h7b, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h8f, 8'h8c, 8'h8c, 8'h8c, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h23, 8'h8e, 8'h81, 8'he, 8'h2b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h63, 8'h0, 8'h16, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h9, 8'h1a, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h2a, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h24, 8'h9a, 8'h9b, 8'h9b, 8'h34, 8'h0, 8'h49, 8'h42, 8'h0, 8'h28, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h23, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h1f, 8'h0, 8'h56, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h22, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h33, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1e, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h76, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h21, 8'h40, 8'h0, 8'h7, 8'h84, 8'h9b, 8'h9b, 8'h77, 8'hb, 8'h0, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h24, 8'h0, 8'h44, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h37, 8'h0, 8'h31, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h1f, 8'h0, 8'h28, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7b, 8'h3, 8'h0, 8'h36, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h78, 8'h1, 8'hb, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h34, 8'h7, 8'h5b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'h7, 8'hb, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h2, 8'h24, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h35, 8'h0, 8'h0, 8'h32, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h20, 8'h93, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h94, 8'h7b, 8'h13, 8'h0, 8'h5f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h20, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h1d, 8'h0, 8'h67, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h29, 8'h0, 8'h0, 8'h3c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h20, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h70, 8'h18, 8'h0, 8'h0, 8'h5b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h93, 8'h91, 8'h91, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h27, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h31, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h17, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h73, 8'h0, 8'h0, 8'h6b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8a, 8'h17, 8'h0, 8'h0, 8'h40, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h96, 8'h93, 8'h92, 8'h96, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h26, 8'h82, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'he, 8'hc, 8'h84, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h5, 8'h25, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h83, 8'hc, 8'h0, 8'h37, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h1f, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h55, 8'h0, 8'h30, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'h2b, 8'h0, 8'h0, 8'h32, 8'h7e, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h24, 8'h0, 8'h1e, 8'h3, 8'h0, 8'h1c, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h40, 8'h0, 8'h1f, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h1e, 8'h0, 8'h5e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2f, 8'h0, 8'h1c, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h1c, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4d, 8'h0, 8'h32, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h42, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h1b, 8'h27, 8'h95, 8'h9b, 8'h40, 8'h0, 8'h37, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h0, 8'h42, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h42, 8'h0, 8'h2f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h93, 8'h95, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h1a, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h10, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h19, 8'h0, 8'h4a, 8'h95, 8'h2d, 8'h0, 8'h0, 8'h15, 8'h85, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h24, 8'hf, 8'h7c, 8'h9a, 8'h76, 8'h2, 8'h21, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h74, 8'h0, 8'h10, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h16, 8'h1c, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h80, 8'h33, 8'h0, 8'h6, 8'h60, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h41, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h89, 8'h82, 8'h87, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h12, 8'h0, 8'h5b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h39, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h26, 8'h0, 8'h0, 8'h69, 8'h99, 8'h79, 8'ha, 8'h0, 8'h18, 8'h85, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h54, 8'h0, 8'h1e, 8'h7e, 8'h4f, 8'h0, 8'h8, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h26, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h25, 8'h0, 8'h44, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h81, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h28, 8'h0, 8'h0, 8'h0, 8'he, 8'h78, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h72, 8'h0, 8'h0, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2f, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8b, 8'h23, 8'h0, 8'h0, 8'h63, 8'h99, 8'h8c, 8'h1c, 8'h0, 8'h0, 8'h61, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h30, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h1c, 8'h0, 8'h67, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6b, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h15, 8'h68, 8'hd, 8'h0, 8'h39, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h44, 8'h0, 8'h2b, 8'h9b, 8'h98, 8'h93, 8'h90, 8'h92, 8'h96, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h3d, 8'h0, 8'h0, 8'h39, 8'h2, 8'h0, 8'h0, 8'h3b, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h41, 8'h0, 8'h22, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2e, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h49, 8'h0, 8'h0, 8'h65, 8'h99, 8'h99, 8'h44, 8'h0, 8'h15, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h71, 8'he, 8'h0, 8'h5a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h4f, 8'h0, 8'h1d, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h1e, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h2d, 8'h0, 8'h40, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h26, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h23, 8'h94, 8'h5c, 8'h0, 8'h0, 8'h0, 8'h37, 8'h84, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h4, 8'h0, 8'h54, 8'h9b, 8'h9a, 8'h35, 8'h0, 8'h0, 8'h19, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h23, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h94, 8'h93, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2c, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h59, 8'h0, 8'h0, 8'h67, 8'h93, 8'h91, 8'h1f, 8'h0, 8'h4f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h4a, 8'h0, 8'h2f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h47, 8'h0, 8'h39, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h1c, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h85, 8'hf, 8'h6, 8'h46, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h85, 8'h98, 8'h9b, 8'h9a, 8'h95, 8'h2a, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h5c, 8'h0, 8'h0, 8'h27, 8'h93, 8'h99, 8'h9a, 8'h9a, 8'h9a, 8'h97, 8'h94, 8'h91, 8'h1d, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h92, 8'h6c, 8'h1f, 8'h0, 8'h35, 8'h7a, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h47, 8'h0, 8'h0, 8'h7, 8'h0, 8'h0, 8'h0, 8'h53, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h79, 8'h0, 8'h17, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h1c, 8'h1a, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h5f, 8'h0, 8'h1c, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h76, 8'h0, 8'h0, 8'h64, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h34, 8'h9b, 8'h7f, 8'h1e, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h8d, 8'h90, 8'h38, 8'h0, 8'h0, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h0, 8'h12, 8'h69, 8'h76, 8'h77, 8'h71, 8'h42, 8'ha, 8'h0, 8'h0, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h52, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h23, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h1f, 8'h95, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2b, 8'h0, 8'h2b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h0, 8'h3a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h79, 8'h59, 8'h5d, 8'h7a, 8'h91, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h22, 8'h0, 8'h68, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h15, 8'h0, 8'h5c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h72, 8'ha, 8'h0, 8'h53, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h84, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h45, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h63, 8'h0, 8'h0, 8'h62, 8'h9b, 8'h9b, 8'h8f, 8'h28, 8'h0, 8'h31, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h5f, 8'h0, 8'hd, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h72, 8'h69, 8'h7e, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h11, 8'h4, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h16, 8'h26, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h92, 8'h9b, 8'h9b, 8'h60, 8'h0, 8'h2b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h14, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'h29, 8'h0, 8'h0, 8'h37, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h4d, 8'ha, 8'h0, 8'h0, 8'h4, 8'h35, 8'h6a, 8'h7f, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6e, 8'h0, 8'h0, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h18, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h66, 8'h0, 8'h8, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h37, 8'h0, 8'h25, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h2c, 8'h0, 8'h4b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1b, 8'h90, 8'h9b, 8'h37, 8'h0, 8'h3b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h14, 8'h0, 8'h5a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h1c, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h30, 8'h0, 8'h35, 8'h9a, 8'h9b, 8'h9a, 8'h61, 8'h0, 8'h4, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h1b, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'he, 8'h29, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1d, 8'h0, 8'h21, 8'h99, 8'h83, 8'h9, 8'h0, 8'h0, 8'h29, 8'h97, 8'h2c, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h15, 8'h0, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h6e, 8'h0, 8'h15, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h5, 8'h79, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h1, 8'h75, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h43, 8'h0, 8'h21, 8'h97, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h0, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h1b, 8'h0, 8'h22, 8'h98, 8'h9b, 8'h68, 8'h0, 8'h0, 8'h0, 8'h58, 8'h29, 8'h0, 8'h42, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h21, 8'h0, 8'h22, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h2b, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h27, 8'h8a, 8'h90, 8'h49, 8'h0, 8'h1, 8'h78, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h1e, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'ha, 8'h28, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h8e, 8'he, 8'h0, 8'h24, 8'h99, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h0, 8'h2b, 8'h29, 8'h0, 8'h3e, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h55, 8'h0, 8'h0, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'hc, 8'h0, 8'h3b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h8c, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h45, 8'h0, 8'h1f, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h27, 8'h0, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h96, 8'h79, 8'h6, 8'h0, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9b, 8'h42, 8'h0, 8'h0, 8'h2a, 8'h38, 8'h0, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h1c, 8'h0, 8'h37, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h8f, 8'h91, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'hd, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6c, 8'h44, 8'h46, 8'h33, 8'h56, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h1f, 8'h0, 8'h5d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hc, 8'h27, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h17, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h95, 8'h9b, 8'h9b, 8'h98, 8'h35, 8'h0, 8'h0, 8'h30, 8'h98, 8'h26, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h40, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8c, 8'h19, 8'h0, 8'h0, 8'h43, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h18, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h48, 8'h0, 8'h1f, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h29, 8'h0, 8'h55, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h0, 8'h6d, 8'h99, 8'h38, 8'h0, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h2d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h19, 8'h0, 8'h0, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h68, 8'h0, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1e, 8'h0, 8'h60, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h12, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2f, 8'h0, 8'h0, 8'h24, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h1a, 8'h0, 8'h0, 8'h30, 8'h9b, 8'h87, 8'h10, 8'h0, 8'h4b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h66, 8'h0, 8'h18, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h20, 8'h9b, 8'h61, 8'h0, 8'h36, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h97, 8'h93, 8'h1b, 8'h0, 8'h1e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h43, 8'h0, 8'h20, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h4d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h1a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7b, 8'h0, 8'h0, 8'h15, 8'h8a, 8'h9b, 8'h5d, 8'h0, 8'h2a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h1b, 8'hc, 8'h7f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h1b, 8'h0, 8'h39, 8'h9b, 8'h93, 8'h24, 8'h23, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h66, 8'h49, 8'hf, 8'h0, 8'h0, 8'h3d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1c, 8'h0, 8'h6d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h93, 8'h1a, 8'h25, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h1d, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h72, 8'h0, 8'h0, 8'h58, 8'h9a, 8'h9b, 8'h61, 8'h0, 8'h31, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h18, 8'hc, 8'h82, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h78, 8'h0, 8'h0, 8'h7a, 8'h9b, 8'h9b, 8'h2d, 8'h0, 8'h63, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h38, 8'h0, 8'h23, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3a, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h9, 8'h0, 8'h5d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h56, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9b, 8'h66, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h1a, 8'hd, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h8f, 8'h8c, 8'h8d, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h37, 8'h0, 8'h1d, 8'h98, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h36, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5b, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h5c, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h14, 8'h2, 8'h7c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h1f, 8'h1d, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9a, 8'h69, 8'h0, 8'h1b, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8d, 8'h10, 8'h0, 8'h1c, 8'h97, 8'h9b, 8'h9b, 8'h67, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h19, 8'hb, 8'h80, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h41, 8'h0, 8'h0, 8'h0, 8'h35, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h20, 8'h0, 8'h20, 8'h9a, 8'h9b, 8'h9b, 8'h7c, 8'h7, 8'h18, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h23, 8'h0, 8'h1e, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h0, 8'h29, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h52, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h22, 8'h0, 8'h25, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h95, 8'h80, 8'h7, 8'h0, 8'h0, 8'h4d, 8'h9b, 8'h9b, 8'h9b, 8'h68, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h15, 8'hd, 8'h81, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h32, 8'h0, 8'h0, 8'h43, 8'h1, 8'h0, 8'h46, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h95, 8'h95, 8'h95, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h1b, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h24, 8'h0, 8'h58, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h11, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h0, 8'h12, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h23, 8'h9, 8'h7e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h78, 8'h0, 8'h0, 8'h42, 8'h98, 8'h94, 8'h91, 8'h84, 8'h1a, 8'h0, 8'h0, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h60, 8'h0, 8'h36, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h68, 8'h0, 8'h1f, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h4a, 8'h0, 8'h1d, 8'h89, 8'h9b, 8'h25, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h88, 8'h44, 8'h11, 8'h19, 8'h17, 8'h3f, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'h2, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2b, 8'h0, 8'h36, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h7, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h21, 8'h0, 8'h39, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h7, 8'h29, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h29, 8'h0, 8'hf, 8'h7c, 8'h5b, 8'hc, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h52, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h52, 8'h0, 8'h29, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'ha, 8'h0, 8'h6c, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h19, 8'h8d, 8'h96, 8'h87, 8'h35, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h22, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h53, 8'h0, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h25, 8'h97, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h0, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h58, 8'h0, 8'h1d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h44, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h21, 8'h16, 8'h87, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h63, 8'h0, 8'h1d, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h26, 8'h0, 8'h46, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h49, 8'h34, 8'h0, 8'h0, 8'h3, 8'h6a, 8'h9a, 8'h9b, 8'h9a, 8'h28, 8'h0, 8'h52, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h0, 8'h1b, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'he, 8'h0, 8'h58, 8'h99, 8'h9b, 8'h3a, 8'h0, 8'h16, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h1c, 8'h0, 8'h63, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h1a, 8'h25, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2b, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h63, 8'h0, 8'h22, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h1b, 8'h0, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h47, 8'h0, 8'h29, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h22, 8'h0, 8'h0, 8'h0, 8'h2, 8'h68, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2d, 8'h0, 8'h3e, 8'h9a, 8'h97, 8'h7b, 8'h61, 8'h72, 8'h8f, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'hc, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3d, 8'h0, 8'h13, 8'h88, 8'h96, 8'h1a, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h47, 8'h0, 8'h37, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h26, 8'h0, 8'h0, 8'h0, 8'hb, 8'h7a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h40, 8'h0, 8'h0, 8'h37, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h31, 8'h0, 8'h35, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h23, 8'h0, 8'h60, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7e, 8'h11, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h29, 8'h0, 8'h33, 8'h96, 8'h33, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h62, 8'h8b, 8'h8f, 8'h95, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h13, 8'h0, 8'h0, 8'h61, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h27, 8'h0, 8'h24, 8'h4d, 8'h0, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8a, 8'hc, 8'h12, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'hd, 8'h82, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h78, 8'h34, 8'h46, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h89, 8'h15, 8'h0, 8'h0, 8'h2a, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h6, 8'h1b, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h2c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h30, 8'h3b, 8'h0, 8'h33, 8'h94, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h70, 8'h91, 8'h92, 8'h93, 8'h99, 8'h9a, 8'h99, 8'h9b, 8'h9b, 8'h98, 8'h8a, 8'h11, 8'h0, 8'h0, 8'h35, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h79, 8'h3, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h21, 8'h0, 8'h3f, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hb, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h16, 8'h0, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2c, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h22, 8'h0, 8'h68, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h40, 8'h0, 8'h0, 8'h0, 8'h21, 8'h91, 8'h9a, 8'h9a, 8'h9b, 8'h8b, 8'h54, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h4d, 8'h7c, 8'h82, 8'h86, 8'h83, 8'h56, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h47, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h4e, 8'h0, 8'h1f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h31, 8'h0, 8'h49, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'he, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h55, 8'h0, 8'h28, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h2a, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h23, 8'h0, 8'h0, 8'h5d, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h18, 8'h0, 8'h79, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h20, 8'h1f, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h52, 8'h0, 8'h0, 8'h75, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h1e, 8'h2a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h24, 8'h0, 8'h4b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h95, 8'h8a, 8'h87, 8'h8d, 8'h92, 8'h95, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h71, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h61, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h13, 8'h26, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5e, 8'h0, 8'h29, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h67, 8'h0, 8'h1d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h58, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h43, 8'h0, 8'h3a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h39, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h1f, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h1b, 8'h0, 8'h69, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h1f, 8'h23, 8'h99, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h6f, 8'h4, 8'h17, 8'h81, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h56, 8'h0, 8'he, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h31, 8'h0, 8'h32, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6d, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h97, 8'h74, 8'hc, 8'h0, 8'h66, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h44, 8'h0, 8'h1, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h98, 8'h3e, 8'h0, 8'h18, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h1e, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h99, 8'h40, 8'h0, 8'h0, 8'h65, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h2e, 8'h0, 8'h6, 8'h73, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h58, 8'h0, 8'hb, 8'h7b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h1b, 8'h0, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h20, 8'h20, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h1f, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h74, 8'h13, 8'h0, 8'h21, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h5d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h91, 8'h8f, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h26, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h7e, 8'h9, 8'h29, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h34, 8'h0, 8'h46, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h85, 8'h2b, 8'h0, 8'h0, 8'h1f, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2d, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h23, 8'h0, 8'h0, 8'h0, 8'h50, 8'h98, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h1f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h35, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h27, 8'hb, 8'h7b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h7a, 8'hb, 8'h0, 8'he, 8'h75, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h83, 8'he, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h53, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h18, 8'h3, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h17, 8'h8c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h1d, 8'h2a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h9a, 8'h95, 8'h55, 8'h0, 8'h0, 8'h45, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h37, 8'h0, 8'h30, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h23, 8'h0, 8'h28, 8'h92, 8'h1e, 8'h0, 8'h16, 8'h8a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h0, 8'h39, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h90, 8'h18, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h91, 8'h1e, 8'h2c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h94, 8'h87, 8'h7c, 8'h7a, 8'h85, 8'h37, 8'h0, 8'h0, 8'h46, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h2, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h93, 8'h90, 8'h8f, 8'h8f, 8'h90, 8'h94, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h0, 8'h2a, 8'h9b, 8'h5e, 8'h0, 8'h0, 8'h1f, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h48, 8'h0, 8'h22, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h54, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h20, 8'h2b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'h12, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h62, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h18, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h8b, 8'h55, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h75, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h22, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h0, 8'h23, 8'h8f, 8'h96, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'hc, 8'h18, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h69, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h1f, 8'h28, 8'h98, 8'h9b, 8'h9b, 8'h99, 8'h95, 8'h68, 8'h0, 8'h0, 8'h2a, 8'h7e, 8'h68, 8'h22, 8'h26, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h93, 8'h8f, 8'h8f, 8'h90, 8'h8f, 8'h90, 8'h8b, 8'h1e, 8'h0, 8'h1e, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h93, 8'h68, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h75, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h21, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9a, 8'h3b, 8'h0, 8'h0, 8'h6, 8'h2e, 8'h54, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h1e, 8'h0, 8'h5e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h20, 8'h22, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h94, 8'h21, 8'h1b, 8'h8c, 8'h9b, 8'h98, 8'h7b, 8'h1b, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h84, 8'h3b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1c, 8'h88, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h86, 8'h41, 8'h0, 8'h0, 8'h0, 8'h9, 8'h46, 8'h80, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h2f, 8'h0, 8'h23, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h25, 8'h0, 8'h29, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h10, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h89, 8'h13, 8'h29, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h34, 8'h0, 8'h38, 8'h92, 8'h50, 8'h0, 8'h0, 8'h1f, 8'h7e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h13, 8'h30, 8'h1c, 8'h0, 8'h0, 8'h0, 8'h29, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h77, 8'h18, 8'h0, 8'h0, 8'h0, 8'h48, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h86, 8'h12, 8'h0, 8'h39, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h0, 8'h19, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h75, 8'h13, 8'h0, 8'h0, 8'h2e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h60, 8'h0, 8'h20, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h4a, 8'h0, 8'h3a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h7f, 8'hc, 8'h0, 8'h0, 8'h0, 8'h0, 8'h63, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h4f, 8'h0, 8'h14, 8'h7b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h90, 8'h33, 8'h0, 8'h0, 8'h3a, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h48, 8'h0, 8'h23, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5e, 8'h0, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h47, 8'h0, 8'h0, 8'h5b, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h15, 8'h13, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h26, 8'h0, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h4d, 8'h0, 8'h0, 8'h31, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h83, 8'h16, 8'h16, 8'h83, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h93, 8'h93, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h93, 8'h91, 8'h60, 8'h0, 8'h0, 8'h2d, 8'h8d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3e, 8'h0, 8'h24, 8'h99, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h1f, 8'h0, 8'h1d, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h96, 8'h26, 8'h0, 8'h0, 8'h60, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h1e, 8'h0, 8'h54, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h21, 8'h24, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h67, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h87, 8'h3b, 8'h0, 8'h0, 8'h45, 8'h90, 8'h97, 8'h9a, 8'h98, 8'h95, 8'h94, 8'h94, 8'h94, 8'h93, 8'h92, 8'h85, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h60, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h3a, 8'h0, 8'h22, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h55, 8'h0, 8'h0, 8'h24, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h1e, 8'h0, 8'h17, 8'h8c, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2b, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h14, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h72, 8'h3, 8'h0, 8'h63, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h71, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h7c, 8'h68, 8'h31, 8'h12, 8'h14, 8'h8, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h20, 8'h72, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h25, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h48, 8'h0, 8'h0, 8'h49, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h6d, 8'h0, 8'h0, 8'h28, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h59, 8'h0, 8'h21, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h57, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h98, 8'h8a, 8'h1f, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h25, 8'h0, 8'h17, 8'h89, 8'h6b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2f, 8'h86, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h20, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h2b, 8'h0, 8'h0, 8'h6c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3e, 8'h0, 8'h0, 8'h4f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h10, 8'h1a, 8'h94, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2c, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h8d, 8'h7b, 8'h5a, 8'h3, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h78, 8'h1, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h99, 8'h4f, 8'h0, 8'h0, 8'h0, 8'h3d, 8'h8a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h11, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8a, 8'h18, 8'h0, 8'h16, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h25, 8'h0, 8'hd, 8'h83, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1c, 8'h0, 8'h6d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h24, 8'h1a, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h95, 8'h8d, 8'h3a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2d, 8'h0, 8'h1a, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8b, 8'h13, 8'h0, 8'h4d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h76, 8'h0, 8'h0, 8'h22, 8'h8f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h68, 8'h0, 8'h0, 8'h24, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h39, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h82, 8'h18, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h40, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h68, 8'h0, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h22, 8'h0, 8'h26, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h0, 8'h18, 8'h8c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h0, 8'h35, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h25, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h82, 8'hd, 8'h29, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h63, 8'h0, 8'h0, 8'h0, 8'hb, 8'h72, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h92, 8'h3e, 8'h0, 8'h0, 8'h14, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h48, 8'h0, 8'h0, 8'h5e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h62, 8'h0, 8'h0, 8'h29, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h2a, 8'h0, 8'h0, 8'h3d, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h69, 8'h0, 8'h20, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h7c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h35, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h61, 8'h0, 8'h0, 8'h1a, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h87, 8'h14, 8'h0, 8'h0, 8'h21, 8'h8b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h24, 8'h0, 8'h1e, 8'h91, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h55, 8'h0, 8'h0, 8'h6b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h1e, 8'h0, 8'h0, 8'h42, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h92, 8'h13, 8'h18, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h5c, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2f, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h59, 8'h0, 8'h0, 8'h16, 8'h85, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h58, 8'h0, 8'h0, 8'h0, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8c, 8'h87, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'h1, 8'h0, 8'h2f, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h22, 8'h0, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h8d, 8'h1c, 8'h0, 8'h0, 8'h36, 8'h8d, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1c, 8'h0, 8'h72, 8'h9b, 8'h9b, 8'h9a, 8'h52, 8'h50, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h14, 8'h89, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6c, 8'h0, 8'h0, 8'h2a, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h73, 8'h2, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h67, 8'h0, 8'h0, 8'h0, 8'h70, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h42, 8'h0, 8'h0, 8'h35, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'ha, 8'h0, 8'h0, 8'h0, 8'h6c, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h20, 8'h0, 8'h49, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h32, 8'h74, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h24, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h1f, 8'h0, 8'h1f, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6f, 8'h0, 8'h0, 8'h0, 8'h39, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h18, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h36, 8'h0, 8'h0, 8'h35, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h99, 8'h99, 8'h97, 8'h2c, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h30, 8'h0, 8'h0, 8'h0, 8'h2d, 8'h8e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h0, 8'h2a, 8'h9a, 8'h9b, 8'h9a, 8'h7b, 8'h31, 8'h52, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h1d, 8'h26, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h93, 8'h26, 8'h0, 8'h0, 8'h5a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h91, 8'h38, 8'h0, 8'h0, 8'h19, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3e, 8'h0, 8'h4d, 8'h33, 8'h0, 8'h23, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h0, 8'h3f, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h7a, 8'h65, 8'h67, 8'h46, 8'h0, 8'h0, 8'h42, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h63, 8'h0, 8'h0, 8'h0, 8'h30, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h4b, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h34, 8'h40, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h7, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h84, 8'h10, 8'h0, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h84, 8'hf, 8'h0, 8'h0, 8'h2b, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h18, 8'h83, 8'h67, 8'h0, 8'h0, 8'h6b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h60, 8'h0, 8'h0, 8'h4d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h90, 8'h1b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'he, 8'h0, 8'h23, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h77, 8'h0, 8'h20, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3a, 8'h3c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4f, 8'h0, 8'h36, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h90, 8'h8a, 8'h8c, 8'h8b, 8'h8f, 8'h94, 8'h95, 8'h96, 8'h95, 8'h74, 8'h2, 8'h0, 8'h0, 8'h66, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h6a, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2d, 8'h17, 8'h82, 8'h9a, 8'h21, 8'h0, 8'h42, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h4e, 8'h0, 8'h0, 8'h66, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h27, 8'h0, 8'h0, 8'h27, 8'h44, 8'h46, 8'h69, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h1d, 8'h0, 8'h21, 8'h95, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h16, 8'h1a, 8'h95, 8'h9b, 8'h9b, 8'h9a, 8'h33, 8'h30, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h34, 8'h0, 8'h51, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h28, 8'h29, 8'h13, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h32, 8'h0, 8'h0, 8'h18, 8'h86, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h5c, 8'h9b, 8'h26, 8'h0, 8'h4a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h43, 8'h0, 8'h0, 8'h5e, 8'h9a, 8'h9b, 8'h9a, 8'h82, 8'h8, 8'h0, 8'h4e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h19, 8'h0, 8'h1f, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1b, 8'h0, 8'h7a, 8'h9b, 8'h9b, 8'h9a, 8'h3b, 8'h26, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h26, 8'h2, 8'h76, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h29, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h94, 8'h77, 8'h7, 8'h0, 8'h0, 8'h34, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3e, 8'h0, 8'h40, 8'h9b, 8'h26, 8'h0, 8'h4b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h54, 8'h0, 8'h10, 8'h80, 8'h9a, 8'h9b, 8'h7a, 8'h2, 8'h4, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7b, 8'h2, 8'h0, 8'h29, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1d, 8'h0, 8'h58, 8'h9a, 8'h9b, 8'h9b, 8'h44, 8'hb, 8'h62, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h21, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7f, 8'hd, 8'h0, 8'h0, 8'h5, 8'h5c, 8'h66, 8'h64, 8'h61, 8'h6d, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h84, 8'h15, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h3c, 8'h0, 8'h38, 8'h9a, 8'h26, 8'h0, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h38, 8'h0, 8'h37, 8'h9b, 8'h9a, 8'h7b, 8'h3, 8'h4, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6a, 8'h0, 8'h0, 8'h31, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h22, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h59, 8'h1, 8'h44, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h31, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h88, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h99, 8'h99, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h93, 8'h4d, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h65, 8'h0, 8'h1e, 8'h80, 8'h16, 8'h0, 8'h6c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h57, 8'h0, 8'h36, 8'h9b, 8'h9b, 8'h80, 8'h8, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h52, 8'h0, 8'h0, 8'h39, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'h15, 8'h3b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h23, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h8f, 8'h31, 8'h0, 8'h0, 8'h0, 8'h66, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h90, 8'h8a, 8'h79, 8'h6c, 8'h6b, 8'h6a, 8'h6c, 8'h79, 8'h8a, 8'h8f, 8'h8e, 8'h60, 8'h0, 8'h0, 8'h0, 8'h15, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h0, 8'h0, 8'h0, 8'h21, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h53, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h92, 8'h91, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h41, 8'h0, 8'h24, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h1e, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h1e, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h62, 8'h0, 8'h0, 8'h0, 8'h1a, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h93, 8'h87, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h20, 8'h0, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h50, 8'h0, 8'h32, 8'h9a, 8'h9b, 8'h9a, 8'h22, 8'h0, 8'h36, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h34, 8'h0, 8'h0, 8'h5d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h99, 8'h4b, 8'h0, 8'h0, 8'h49, 8'h8f, 8'h97, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h60, 8'h0, 8'h21, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h25, 8'h2c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h7d, 8'hc, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h91, 8'h5d, 8'h1, 8'h0, 8'h2f, 8'h90, 8'h95, 8'h96, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h92, 8'h91, 8'h84, 8'h51, 8'h2, 8'h0, 8'h0, 8'h0, 8'h0, 8'h12, 8'h55, 8'h78, 8'h75, 8'h76, 8'h77, 8'h3a, 8'h0, 8'h0, 8'h0, 8'hd, 8'h6c, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h5, 8'h60, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4d, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h0, 8'h0, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4c, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7c, 8'h0, 8'h20, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h27, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h60, 8'h0, 8'h36, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h0, 8'h26, 8'h36, 8'h5b, 8'h96, 8'h98, 8'h98, 8'h95, 8'h91, 8'h74, 8'h26, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h5d, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h2c, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h53, 8'h0, 8'h0, 8'h32, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h23, 8'h0, 8'h12, 8'h76, 8'h24, 8'h0, 8'h0, 8'h0, 8'h70, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h11, 8'h1c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h2d, 8'h1d, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h47, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h91, 8'h92, 8'h35, 8'h0, 8'h28, 8'h60, 8'h4f, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2, 8'h55, 8'h8c, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h97, 8'h98, 8'h96, 8'h98, 8'h97, 8'h96, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h76, 8'h3, 8'h18, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h63, 8'h0, 8'h1d, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h4, 8'h0, 8'h3, 8'h75, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h8b, 8'h13, 8'h0, 8'h36, 8'h9b, 8'h9b, 8'h87, 8'h16, 8'h0, 8'h0, 8'h49, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h18, 8'h14, 8'h91, 8'h9b, 8'h9a, 8'h9b, 8'h2e, 8'h6, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h58, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h59, 8'h93, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h96, 8'h95, 8'h92, 8'h8f, 8'h8c, 8'h89, 8'h8b, 8'h87, 8'h6b, 8'h4b, 8'h45, 8'h47, 8'h43, 8'h45, 8'h44, 8'h4d, 8'h71, 8'h8d, 8'h93, 8'h96, 8'h96, 8'h98, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h29, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7b, 8'h5, 8'h19, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h30, 8'h0, 8'h0, 8'h6, 8'h75, 8'h97, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h6d, 8'h0, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h31, 8'h0, 8'h0, 8'h3e, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1c, 8'h1, 8'h7c, 8'h9b, 8'h9b, 8'h9b, 8'h3a, 8'h1, 8'h62, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h4, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h93, 8'h8c, 8'h69, 8'h3e, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h2c, 8'h44, 8'h54, 8'h7a, 8'h8f, 8'h92, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h72, 8'h0, 8'h1, 8'h75, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h76, 8'h0, 8'h11, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h22, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h93, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h5, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h35, 8'h0, 8'h0, 8'h4f, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h1c, 8'h0, 8'h6b, 8'h9b, 8'h9b, 8'h9b, 8'h42, 8'h0, 8'h4e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h11, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h8e, 8'h89, 8'h83, 8'h87, 8'h92, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h93, 8'h8d, 8'h7d, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h1e, 8'h1f, 8'h22, 8'h20, 8'h20, 8'h6, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h37, 8'h7e, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h25, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h92, 8'h1a, 8'h0, 8'h6c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h2f, 8'h0, 8'h0, 8'h0, 8'h3a, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h5, 8'h7b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h67, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1d, 8'h0, 8'h5c, 8'h9b, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h26, 8'h1b, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h78, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'hc, 8'h77, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h93, 8'h8f, 8'h81, 8'h44, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h19, 8'h54, 8'h7d, 8'h94, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h89, 8'h5a, 8'h2c, 8'h1d, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h15, 8'h77, 8'h90, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h3e, 8'h0, 8'ha, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h28, 8'h0, 8'h60, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h71, 8'h0, 8'h0, 8'h3, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5f, 8'h0, 8'h4, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h3d, 8'h0, 8'h0, 8'h0, 8'h36, 8'h94, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1f, 8'h0, 8'h49, 8'h9b, 8'h9a, 8'h9b, 8'h63, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h1d, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h83, 8'h88, 8'h80, 8'h28, 8'h9, 8'h4f, 8'h83, 8'h8e, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h67, 8'h93, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h94, 8'h92, 8'h90, 8'h87, 8'h51, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h16, 8'h68, 8'h92, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h5b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h92, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h67, 8'h0, 8'h0, 8'h54, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h4a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h3e, 8'h0, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h1, 8'h78, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h38, 8'h0, 8'h0, 8'h19, 8'h85, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h0, 8'h3c, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h9, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h21, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h42, 8'h0, 8'h2a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h50, 8'h0, 8'h0, 8'h0, 8'h1, 8'h6a, 8'h8e, 8'h91, 8'h96, 8'h98, 8'h94, 8'h92, 8'h92, 8'h92, 8'h91, 8'h92, 8'h90, 8'h87, 8'h66, 8'h21, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h66, 8'h92, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h11, 8'h0, 8'h0, 8'h0, 8'h7, 8'h74, 8'h97, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8e, 8'h16, 8'h0, 8'h2b, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h44, 8'h0, 8'h38, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h79, 8'h1, 8'h0, 8'h23, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h62, 8'h0, 8'h5, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h53, 8'h0, 8'h0, 8'h0, 8'h20, 8'h6e, 8'h88, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h34, 8'h9a, 8'h9b, 8'h9b, 8'h7f, 8'h13, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h25, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h47, 8'h0, 8'h0, 8'h42, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h4a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h4e, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h95, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h93, 8'h34, 8'h0, 8'h0, 8'h0, 8'h40, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h34, 8'h0, 8'ha, 8'h7f, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5f, 8'h0, 8'h2f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h1d, 8'h0, 8'he, 8'h83, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h6a, 8'h0, 8'h10, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h73, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h92, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9a, 8'h88, 8'h1a, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h25, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h1b, 8'h0, 8'h1b, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h43, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3c, 8'h74, 8'h8e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7c, 8'he, 8'h0, 8'h0, 8'h12, 8'h84, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h20, 8'h0, 8'h31, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h21, 8'h1e, 8'h8e, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2f, 8'h0, 8'h0, 8'h5d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h6b, 8'h0, 8'hf, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h67, 8'h11, 8'h0, 8'h0, 8'h0, 8'h2e, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2d, 8'h0, 8'h29, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h20, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h24, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6b, 8'h0, 8'h0, 8'h31, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h73, 8'h39, 8'h28, 8'h5d, 8'h80, 8'h7f, 8'h83, 8'h82, 8'h80, 8'h8d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h4c, 8'h0, 8'h0, 8'h23, 8'h94, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h75, 8'h0, 8'h0, 8'h63, 8'h9b, 8'h95, 8'h92, 8'h90, 8'h91, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'hf, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h54, 8'h0, 8'h0, 8'h37, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h66, 8'h0, 8'h8, 8'h7e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h2b, 8'h0, 8'h9, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h32, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h26, 8'h2f, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h25, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h26, 8'h0, 8'h5, 8'h83, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h0, 8'h3b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h39, 8'h0, 8'h16, 8'h86, 8'h88, 8'h31, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h91, 8'h9a, 8'h9b, 8'h9b, 8'h29, 8'h11, 8'h7f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7c, 8'h4, 8'h0, 8'h22, 8'h94, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h62, 8'h0, 8'hb, 8'h80, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h46, 8'h0, 8'h5, 8'h7a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h37, 8'h0, 8'h25, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h27, 8'h2b, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h5, 8'h0, 8'h20, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h15, 8'h8a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h0, 8'h0, 8'he, 8'h7e, 8'h9b, 8'h9b, 8'h2a, 8'hf, 8'h7d, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h25, 8'h0, 8'h0, 8'h5c, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h5d, 8'h0, 8'h7, 8'h7e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3c, 8'h0, 8'h2, 8'h79, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h40, 8'h0, 8'h24, 8'h9a, 8'h9b, 8'h9a, 8'h97, 8'h25, 8'h27, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h57, 8'h0, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h70, 8'h0, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h0, 8'h0, 8'h18, 8'h81, 8'h9b, 8'h9b, 8'h9a, 8'h43, 8'h0, 8'h2a, 8'h97, 8'h9b, 8'h2a, 8'hf, 8'h7d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h65, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h96, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h3b, 8'h0, 8'h13, 8'h89, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h17, 8'h0, 8'h17, 8'h8a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h25, 8'h20, 8'h90, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h26, 8'h0, 8'h0, 8'h6d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h88, 8'h73, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h28, 8'h0, 8'h4c, 8'h99, 8'h2a, 8'h5, 8'h72, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h35, 8'h8d, 8'h99, 8'h99, 8'h9b, 8'h99, 8'h26, 8'h0, 8'h25, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h4e, 8'h0, 8'h0, 8'h3f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h3f, 8'h0, 8'h24, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h27, 8'h22, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h89, 8'ha, 8'h0, 8'h1d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h0, 8'h29, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7d, 8'hb, 8'h22, 8'h7e, 8'h17, 8'h19, 8'h89, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h52, 8'h0, 8'h0, 8'h0, 8'h0, 8'h58, 8'h72, 8'h78, 8'h5e, 8'h0, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h93, 8'h1e, 8'h0, 8'h11, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h28, 8'h1d, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h5d, 8'h0, 8'h0, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h0, 8'h1c, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h32, 8'h0, 8'h0, 8'h0, 8'h3b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7d, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h8, 8'h7a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h66, 8'h0, 8'h0, 8'h31, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3e, 8'h0, 8'h23, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h18, 8'h88, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h99, 8'h2f, 8'h0, 8'h0, 8'h52, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3a, 8'h0, 8'h18, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h29, 8'h0, 8'h20, 8'h86, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h41, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1, 8'h6b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4f, 8'h0, 8'h0, 8'h60, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h40, 8'h0, 8'h25, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h18, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h21, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h90, 8'h8f, 8'h90, 8'h93, 8'h97, 8'h9a, 8'h9b, 8'h9a, 8'h9a, 8'h97, 8'h1d, 8'h0, 8'h0, 8'h7c, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3d, 8'h0, 8'h14, 8'h8b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h98, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4b, 8'h0, 8'h0, 8'h5c, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h3a, 8'h0, 8'h24, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h18, 8'h88, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h25, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h94, 8'h29, 8'h0, 8'h0, 8'h0, 8'h0, 8'h42, 8'h84, 8'h93, 8'h99, 8'h9b, 8'h8b, 8'h10, 8'h0, 8'h14, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2f, 8'h0, 8'h1c, 8'h90, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h56, 8'h0, 8'h0, 8'h2a, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h37, 8'h0, 8'h26, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h1a, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h21, 8'h24, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8f, 8'h74, 8'h5d, 8'h47, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h65, 8'h95, 8'h6e, 8'h0, 8'h0, 8'h20, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h14, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h18, 8'h0, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h0, 8'h28, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h1a, 8'h89, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h25, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h79, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h0, 8'h0, 8'h0, 8'h25, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h62, 8'h0, 8'h0, 8'h51, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h42, 8'h0, 8'h0, 8'h12, 8'h80, 8'h93, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h93, 8'h90, 8'h92, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2b, 8'h0, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h28, 8'h22, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h24, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h18, 8'h8d, 8'h9a, 8'h9a, 8'h7b, 8'hb, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h46, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h12, 8'h87, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h94, 8'h26, 8'h0, 8'h0, 8'h0, 8'h6, 8'h54, 8'h80, 8'h8c, 8'h8e, 8'h92, 8'h96, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h89, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h4e, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h28, 8'h0, 8'h30, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h26, 8'h23, 8'h92, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h22, 8'h22, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h27, 8'h0, 8'h0, 8'h0, 8'h0, 8'h27, 8'h81, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h97, 8'h39, 8'h0, 8'h0, 8'h0, 8'h0, 8'h1d, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h26, 8'h0, 8'h28, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h85, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h31, 8'h74, 8'h8b, 8'h91, 8'h94, 8'h98, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h86, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h6a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9a, 8'h22, 8'h0, 8'h36, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h24, 8'h23, 8'h93, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h1c, 8'h91, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h5c, 8'h0, 8'h0, 8'hd, 8'h88, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h5c, 8'h5, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h0, 8'h29, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h7a, 8'h2a, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h4f, 8'h79, 8'h8b, 8'h98, 8'h9a, 8'h98, 8'h3e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h14, 8'h38, 8'h0, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1f, 8'h0, 8'h42, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h23, 8'h28, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h11, 8'h84, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h90, 8'h11, 8'h0, 8'h1, 8'h7e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h25, 8'h0, 8'h24, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8d, 8'h73, 8'h64, 8'h3f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h52, 8'h96, 8'h53, 8'h0, 8'h0, 8'h0, 8'h1f, 8'h7d, 8'h9b, 8'h92, 8'h19, 8'h0, 8'h2c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1e, 8'h0, 8'h4f, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h1f, 8'h2a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h28, 8'h1, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h28, 8'h0, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h0, 8'h0, 8'h45, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h95, 8'h87, 8'h6d, 8'h48, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h39, 8'h0, 8'h0, 8'h11, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h20, 8'h0, 8'h2a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1d, 8'h0, 8'h65, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h19, 8'h2c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h30, 8'h0, 8'h5f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h18, 8'h0, 8'h14, 8'h90, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h1f, 8'h0, 8'h2a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h74, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h67, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h21, 8'h0, 8'h24, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1b, 8'h0, 8'h78, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h10, 8'h2d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3a, 8'h0, 8'h44, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2b, 8'h0, 8'h0, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h23, 8'h0, 8'h2c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h35, 8'h0, 8'h0, 8'h60, 8'h90, 8'h90, 8'h90, 8'h92, 8'h96, 8'h97, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h1a, 8'hf, 8'h8b, 8'h9b, 8'h9a, 8'h9b, 8'h74, 8'h5, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h55, 8'h0, 8'h39, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h0, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7f, 8'ha, 8'h0, 8'h38, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h87, 8'h77, 8'h89, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h7c, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h28, 8'h48, 8'h6f, 8'h87, 8'h90, 8'h96, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h17, 8'h1b, 8'h96, 8'h9b, 8'h9b, 8'h9b, 8'h69, 8'h0, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h6d, 8'h0, 8'h2d, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h59, 8'h0, 8'h0, 8'h29, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h2b, 8'h0, 8'h8, 8'h7d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h5f, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h34, 8'h86, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h84, 8'h5, 8'h1e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h59, 8'h0, 8'h37, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8c, 8'h18, 8'h2b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h37, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h65, 8'h0, 8'h0, 8'h39, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h8e, 8'h88, 8'h88, 8'h7d, 8'h56, 8'h36, 8'h8, 8'h0, 8'h0, 8'h0, 8'h0, 8'h25, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6b, 8'h0, 8'h21, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h46, 8'h0, 8'h3d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h97, 8'h20, 8'h28, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h99, 8'h33, 8'h0, 8'h0, 8'h4e, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h91, 8'h1c, 8'h0, 8'h23, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h70, 8'h0, 8'h0, 8'h23, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h4a, 8'h0, 8'h22, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h3c, 8'h0, 8'h4b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h24, 8'h28, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h77, 8'h0, 8'h0, 8'h14, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h90, 8'h1d, 8'h0, 8'h0, 8'h4f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h70, 8'h0, 8'h0, 8'h0, 8'h66, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h0, 8'h27, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h27, 8'h28, 8'h99, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h30, 8'h0, 8'h0, 8'h34, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h90, 8'h1f, 8'h0, 8'h0, 8'h41, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h98, 8'h59, 8'h0, 8'h0, 8'h0, 8'h5d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h24, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h1, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h1f, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h97, 8'h20, 8'h0, 8'h0, 8'h4c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h8c, 8'h19, 8'h0, 8'h0, 8'h44, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h58, 8'h0, 8'h0, 8'h0, 8'h6f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1f, 8'h0, 8'h4d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h13, 8'h82, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h9, 8'h6e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h21, 8'h0, 8'h0, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h2e, 8'h0, 8'h0, 8'h3d, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h1b, 8'h0, 8'h1, 8'h75, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h1c, 8'h0, 8'h72, 8'h9b, 8'h9a, 8'h9b, 8'h96, 8'h25, 8'h22, 8'h90, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4c, 8'h0, 8'h47, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h2f, 8'h0, 8'h0, 8'h2e, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h56, 8'h0, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h56, 8'h0, 8'h0, 8'h45, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h96, 8'h18, 8'h13, 8'h8f, 8'h9b, 8'h9a, 8'h9b, 8'h8c, 8'h1a, 8'h29, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h79, 8'h11, 8'h34, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h76, 8'h0, 8'h0, 8'h0, 8'h3e, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h26, 8'h0, 8'h16, 8'h8c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2b, 8'h0, 8'he, 8'h83, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h2, 8'h1e, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h7a, 8'hb, 8'h2e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h20, 8'h2c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h48, 8'h0, 8'h0, 8'h0, 8'h5b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h2e, 8'h0, 8'h0, 8'h4d, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h91, 8'h1a, 8'h0, 8'h1f, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h5d, 8'h0, 8'h21, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h60, 8'h0, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h26, 8'h29, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h4d, 8'h0, 8'h0, 8'h27, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h14, 8'h0, 8'h1, 8'h77, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h6c, 8'h0, 8'h0, 8'h31, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h35, 8'h0, 8'h26, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h40, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h29, 8'h29, 8'h99, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h97, 8'h1b, 8'h0, 8'h10, 8'h8e, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h72, 8'h0, 8'h0, 8'h52, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h95, 8'h90, 8'h90, 8'h91, 8'h90, 8'h8f, 8'h90, 8'h91, 8'h94, 8'h98, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h38, 8'h0, 8'h0, 8'h53, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h20, 8'h0, 8'h37, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h35, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h33, 8'h1f, 8'h82, 8'h9b, 8'h9b, 8'h9a, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h98, 8'h23, 8'h0, 8'h0, 8'h79, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h72, 8'h0, 8'h0, 8'h5c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hb, 8'h4d, 8'h82, 8'h95, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h20, 8'h0, 8'hf, 8'h82, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h1e, 8'h0, 8'h64, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h2a, 8'h5, 8'h72, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h4d, 8'h1, 8'h50, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h96, 8'h1f, 8'h0, 8'h0, 8'h73, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h74, 8'h0, 8'h0, 8'h59, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3c, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'he, 8'h6b, 8'h92, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8a, 8'h12, 8'h0, 8'h24, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h98, 8'h18, 8'hd, 8'h89, 8'h9b, 8'h9b, 8'h9a, 8'h99, 8'h25, 8'h1b, 8'h8b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h81, 8'h1d, 8'h39, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h92, 8'h1a, 8'h0, 8'h0, 8'h76, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h6e, 8'h0, 8'h0, 8'h57, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h94, 8'h1e, 8'h0, 8'h1e, 8'h8c, 8'h91, 8'h8c, 8'h8b, 8'h7f, 8'h45, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h10, 8'h75, 8'h97, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h77, 8'h0, 8'h0, 8'h2c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h0, 8'h1f, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h8f, 8'h1e, 8'h2c, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h2f, 8'h34, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h5c, 8'h0, 8'h0, 8'h1a, 8'h95, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h64, 8'h0, 8'h0, 8'h61, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h7a, 8'h2, 8'h0, 8'h48, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h80, 8'h28, 8'h0, 8'h0, 8'h0, 8'h0, 8'h45, 8'h8a, 8'h99, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h59, 8'h0, 8'h0, 8'h3a, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h49, 8'h0, 8'h21, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h76, 8'hc, 8'h32, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h31, 8'h34, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h9b, 8'h98, 8'h24, 8'h0, 8'h0, 8'h43, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h56, 8'h0, 8'h1f, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h7a, 8'h2, 8'h0, 8'h60, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h86, 8'h20, 8'h0, 8'h0, 8'h0, 8'h0, 8'h68, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h65, 8'h0, 8'h0, 8'h33, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h27, 8'h0, 8'h2f, 8'h9b, 8'h9a, 8'h9b, 8'h9b, 8'h51, 8'h0, 8'h3e, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h3f, 8'h36, 8'h8f, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h88, 8'h13, 8'h0, 8'h1e, 8'h94, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h99, 8'h8b, 8'h8d, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h86, 8'h14, 8'h0, 8'h70, 8'h9a, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h95, 8'h4e, 8'h0, 8'h0, 8'h0, 8'h0, 8'h56, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h8d, 8'h1c, 8'h0, 8'h2a, 8'h98, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h23, 8'h0, 8'h55, 8'h9b, 8'h9b, 8'h9b, 8'h9a, 8'h3e, 8'h0, 8'h5c, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h9b, 8'h0, 
		8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 
		8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0 

        };

	assign data = ROM[addr];

endmodule