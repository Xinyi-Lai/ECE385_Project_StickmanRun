module digits_rom ( input [7:0] addr, output [7:0] data);

	parameter ROM_LENGTH = 16*10;
	parameter DATA_WIDTH = 8;

	// ROM definition				
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {

		// code x0
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11001110, // 5 **  ***
		8'b11011110, // 6 ** ****
		8'b11110110, // 7 **** **
		8'b11100110, // 8 ***  **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x1
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00011000, // 2
		8'b00111000, // 3
		8'b01111000, // 4    **
		8'b00011000, // 5   ***
		8'b00011000, // 6  ****
		8'b00011000, // 7    **
		8'b00011000, // 8    **
		8'b00011000, // 9    **
		8'b00011000, // a    **
		8'b01111110, // b    **
		8'b00000000, // c    **
		8'b00000000, // d  ******
		8'b00000000, // e
		8'b00000000, // f
		// code x2
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b00000110, // 4      **
		8'b00001100, // 5     **
		8'b00011000, // 6    **
		8'b00110000, // 7   **
		8'b01100000, // 8  **
		8'b11000000, // 9 **
		8'b11000110, // a **   **
		8'b11111110, // b *******
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x3
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b00000110, // 4      **
		8'b00000110, // 5      **
		8'b00111100, // 6   ****
		8'b00000110, // 7      **
		8'b00000110, // 8      **
		8'b00000110, // 9      **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x4
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00001100, // 2     **
		8'b00011100, // 3    ***
		8'b00111100, // 4   ****
		8'b01101100, // 5  ** **
		8'b11001100, // 6 **  **
		8'b11111110, // 7 *******
		8'b00001100, // 8     **
		8'b00001100, // 9     **
		8'b00001100, // a     **
		8'b00011110, // b    ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x5
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111110, // 2 *******
		8'b11000000, // 3 **
		8'b11000000, // 4 **
		8'b11000000, // 5 **
		8'b11111100, // 6 ******
		8'b00000110, // 7      **
		8'b00000110, // 8      **
		8'b00000110, // 9      **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x6
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111000, // 2   ***
		8'b01100000, // 3  **
		8'b11000000, // 4 **
		8'b11000000, // 5 **
		8'b11111100, // 6 ******
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x7
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111110, // 2 *******
		8'b11000110, // 3 **   **
		8'b00000110, // 4      **
		8'b00000110, // 5      **
		8'b00001100, // 6     **
		8'b00011000, // 7    **
		8'b00110000, // 8   **
		8'b00110000, // 9   **
		8'b00110000, // a   **
		8'b00110000, // b   **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x8
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11000110, // 5 **   **
		8'b01111100, // 6  *****
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// code x9
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11000110, // 5 **   **
		8'b01111110, // 6  ******
		8'b00000110, // 7      **
		8'b00000110, // 8      **
		8'b00000110, // 9      **
		8'b00001100, // a     **
		8'b01111000, // b  ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000 // f
	};

	assign data = ROM[addr];

endmodule  




module stickman_rom ( input [9:0] addr, output [55:0] data);

	//parameter ADDR_WIDTH = 10;
	parameter ROM_LENGTH = 80*9;	// 720
	parameter DATA_WIDTH = 56;
				
	// ROM definition: height: 80*9, width: 56
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {
		// height: 80, width: 56
		//Page 1
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000100000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000011100000000000,
		56'b00000000000000000000000000001111111110000111110000000000,
		56'b00000000000000000000000000011111111000000111110000000000,
		56'b00000000000000000000000011111111100000001111110000000000,
		56'b00000000000000000000011111111111100000001111100000000000,
		56'b00000000000000000001111111111111110000011111100000000000,
		56'b00000000000000001111111111111111111000011111000000000000,
		56'b00000000000000001111111111111111111100111111000000000000,
		56'b00000000000000011111111110011111111100111110000000000000,
		56'b00000000000000011111110000011111111111111110000000000000,
		56'b00000000000000011111000000011111111111111100000000000000,
		56'b00000000000000011111000000011111111111111100000000000000,
		56'b00000000000000011111000000011111011111111000000000000000,
		56'b00000000000000011111000000011111001111111000000000000000,
		56'b00000000000000111110000000011110001111110000000000000000,
		56'b00000000000000111110000000011110000111110000000000000000,
		56'b00000000000000111110000000111110000111100000000000000000,
		56'b00000000000000111110000000111110000001000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111100000000111110000000000000000000000000,
		56'b00000000000001111100000000111110000000000000000000000000,
		56'b00000000000001111100000000111110000000000000000000000000,
		56'b00000000000001111100000000111110000000000000000000000000,
		56'b00000000000000111100000001111110000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111111000000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000011111111111111111110000000000000,
		56'b00000000000000000000000011111111111111111111110000000000,
		56'b00000000000000000000000011111001111111111111111000000000,
		56'b00000000000000000000000111111000000111111111111000000000,
		56'b00000000000000000000000111110000000000011111111000000000,
		56'b00000000000000000000001111110000000000001111110000000000,
		56'b00000000000000000000001111100000000000001111100000000000,
		56'b00000000000000000000001111100000000000011111100000000000,
		56'b00000000000000000000011111100000000000111111000000000000,
		56'b00000000000000000000011111000000000000111111000000000000,
		56'b00000000000000000000111111000000000001111110000000000000,
		56'b00000000000000000000111110000000000001111100000000000000,
		56'b00000000000000000000111110000000000011111100000000000000,
		56'b00000000000000000001111100000000000111111000000000000000,
		56'b00000000000000000011111100000000000111110000000000000000,
		56'b00000000000000000111111100000000001111110000000000000000,
		56'b00000000000000011111111000000000011111100000000000000000,
		56'b00000000000000111111110000000000011111100000000000000000,
		56'b00000000000001111111100000000000011111110000000000000000,
		56'b00000000000011111111000000000000011111110000000000000000,
		56'b00000000000111111100000000000000000111110000000000000000,
		56'b00000000011111111000000000000000000011110000000000000000,
		56'b00000000111111110000000000000000000001100000000000000000,
		56'b00000001111111000000000000000000000000000000000000000000,
		56'b00000011111110000000000000000000000000000000000000000000,
		56'b00000111111100000000000000000000000000000000000000000000,
		56'b00000111111000000000000000000000000000000000000000000000,
		56'b00000011111000000000000000000000000000000000000000000000,
		56'b00000011111000000000000000000000000000000000000000000000,
		56'b00000011111000000000000000000000000000000000000000000000,
		56'b00000001111000000000000000000000000000000000000000000000,
		56'b00000000100000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 2
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000011111000000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100111100000000000,
		56'b00000000000000000000000000111111111111101111100000000000,
		56'b00000000000000000000000000111111111111001111100000000000,
		56'b00000000000000000000000000011111111110001111100000000000,
		56'b00000000000000000000000000001111111100001111100000000000,
		56'b00000000000000000000000000011111110000011111000000000000,
		56'b00000000000000000000000011111111110000011111000000000000,
		56'b00000000000000000000001111111111111000011111000000000000,
		56'b00000000000000000001111111111111111100011111000000000000,
		56'b00000000000000000111111111111111111110111111000000000000,
		56'b00000000000000001111111111111111111111111110000000000000,
		56'b00000000000000001111111110011111111111111110000000000000,
		56'b00000000000000001111111000011111011111111110000000000000,
		56'b00000000000000001111000000011111001111111110000000000000,
		56'b00000000000000011111000000011111000111111110000000000000,
		56'b00000000000000011111000000011111000011111100000000000000,
		56'b00000000000000011111000000011110000001111100000000000000,
		56'b00000000000000011111000000011110000000111000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000111111000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000000111110000000000000000000000000,
		56'b00000000000000111110000001111100000000000000000000000000,
		56'b00000000000000011100000001111111100000000000000000000000,
		56'b00000000000000000000000001111111111110000000000000000000,
		56'b00000000000000000000000011111111111111110000000000000000,
		56'b00000000000000000000000011111111111111111111100000000000,
		56'b00000000000000000000000111111111111111111111110000000000,
		56'b00000000000000000000001111110000111111111111111000000000,
		56'b00000000000000000000001111100000000011111111111000000000,
		56'b00000000000000000000011111100000000000001111111000000000,
		56'b00000000000000000000111111000000000000000011111000000000,
		56'b00000000000000000000111110000000000000000111110000000000,
		56'b00000000000000000001111110000000000000000111110000000000,
		56'b00000000000000000011111100000000000000000111110000000000,
		56'b00000000000000000011111100000000000000000111110000000000,
		56'b00000000000000000111111000000000000000000111110000000000,
		56'b00000000000000001111110000000000000000000111110000000000,
		56'b00000000000000011111100000000000000000001111100000000000,
		56'b00000000000001111111100000000000000000001111100000000000,
		56'b00000000000011111111000000000000000000001111100000000000,
		56'b00000000000111111110000000000000000000001111100000000000,
		56'b00000000011111111100000000000000000000001111100000000000,
		56'b00000000111111110000000000000000000000001111100000000000,
		56'b00000011111111100000000000000000000000011111000000000000,
		56'b00000111111110000000000000000000000000011111100000000000,
		56'b00011111111100000000000000000000000000011111110000000000,
		56'b00111111111000000000000000000000000000001111111000000000,
		56'b00111111100000000000000000000000000000000111111000000000,
		56'b00111111000000000000000000000000000000000001110000000000,
		56'b00111110000000000000000000000000000000000000000000000000,
		56'b00111110000000000000000000000000000000000000000000000000,
		56'b00111110000000000000000000000000000000000000000000000000,
		56'b00011110000000000000000000000000000000000000000000000000,
		56'b00001100000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 3
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111000000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111101000000000000000,
		56'b00000000000000000000000001111111111111111100000000000000,
		56'b00000000000000000000000000111111111111111110000000000000,
		56'b00000000000000000000000000111111111111111110000000000000,
		56'b00000000000000000000000000011111111111111110000000000000,
		56'b00000000000000000000000000011111111110111110000000000000,
		56'b00000000000000000000000000001111111100111110000000000000,
		56'b00000000000000000000000000011111110000111110000000000000,
		56'b00000000000000000000000001111111110000111110000000000000,
		56'b00000000000000000000000111111111111000111110000000000000,
		56'b00000000000000000000011111111111111110111110000000000000,
		56'b00000000000000000001111111111111111111111110000000000000,
		56'b00000000000000000011111111111111111111111110000000000000,
		56'b00000000000000001111111111011111011111111110000000000000,
		56'b00000000000000001111111100011111001111111110000000000000,
		56'b00000000000000001111110000011111000111111110000000000000,
		56'b00000000000000001111100000011111000011111110000000000000,
		56'b00000000000000001111100000011111000000111110000000000000,
		56'b00000000000000001111100000011110000000011100000000000000,
		56'b00000000000000000111100000011110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110001111100000000000000000000000000,
		56'b00000000000000000111110001111111100000000000000000000000,
		56'b00000000000000000011100001111111111100000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111111110000000000000,
		56'b00000000000000000000000011111111111111111111100000000000,
		56'b00000000000000000000000011111000011111111111110000000000,
		56'b00000000000000000000000111111000000111111111111000000000,
		56'b00000000000000000000000111110000000000011111111000000000,
		56'b00000000000000000000000111110000000000000011111000000000,
		56'b00000000000000000000001111100000000000000011111000000000,
		56'b00000000000000000000001111100000000000000011111000000000,
		56'b00000000000000000000001111100000000000000011111000000000,
		56'b00000000000000000000011111100000000000000001111000000000,
		56'b00000000000000000000011111000000000000000001111100000000,
		56'b00000000000000000000011111000000000000000001111100000000,
		56'b00000000000000000000111110000000000000000001111100000000,
		56'b00000000000000011111111110000000000000000001111100000000,
		56'b00000000011111111111111110000000000000000001111100000000,
		56'b00001111111111111111111110000000000000000001111100000000,
		56'b00011111111111111111111100000000000000000000111100000000,
		56'b00011111111111111111100000000000000000000000111110000000,
		56'b00111111111111110000000000000000000000000000111110000000,
		56'b00111111000000000000000000000000000000000000111111110000,
		56'b00111110000000000000000000000000000000000000111111110000,
		56'b00111100000000000000000000000000000000000000111111110000,
		56'b00111100000000000000000000000000000000000000011111110000,
		56'b00000000000000000000000000000000000000000000000001000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 4
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000111111111110000000000000000000000,
		56'b00000000000000000000001111111111110000000000000000000000,
		56'b00000000000000000000011111111111110000000000000000000000,
		56'b00000000000000000000111111111111110000000000111000000000,
		56'b00000000000000000000111111011111110000011111111100000000,
		56'b00000000000000000001111110011111111011111111111100000000,
		56'b00000000000000000001111100011111111111111111111100000000,
		56'b00000000000000000001111100111111111111111111111000000000,
		56'b00000000000000000000111100111111111111111111000000000000,
		56'b00000000000000000000111110111111111111110000000000000000,
		56'b00000000000000000000111110111111111100000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111110000000000000000000000000,
		56'b00000000000000000000111110111100000000000000000000000000,
		56'b00000000000000000000011111111100000000000000000000000000,
		56'b00000000000000000000011111111110000000000000000000000000,
		56'b00000000000000000000011111111111000000000000000000000000,
		56'b00000000000000000000011111111111100000000000000000000000,
		56'b00000000000000000000011111111111110000000000000000000000,
		56'b00000000000000000000001111111111111000000000000000000000,
		56'b00000000000000000000000001111111111100000000000000000000,
		56'b00000000000000000000000011111011111110000000000000000000,
		56'b00000000000000000000000011111001111111000000000000000000,
		56'b00000000000000000000000011111000111111110000000000000000,
		56'b00000000000000000000000011111000011111111000000000000000,
		56'b00000000000000000000000011111000000111111100000000000000,
		56'b00000000000000000000000011111000000011111110000000000000,
		56'b00000000000000000000000011110000000001111110000000000000,
		56'b00000011111100000000000111110000000000111110000000000000,
		56'b00000111111111111100000111110000000000011111000000000000,
		56'b00001111111111111111111111110000000000011111000000000000,
		56'b00001111111111111111111111110000000000011111100000000000,
		56'b00011111111111111111111111110000000000001111100000000000,
		56'b00001111000001111111111111100000000000001111110000000000,
		56'b00000110000000000011111111100000000000000111110000000000,
		56'b00000000000000000000000111000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000111111000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000001111100000000,
		56'b00000000000000000000000000000000000000000001111100000000,
		56'b00000000000000000000000000000000000000000001111100000000,
		56'b00000000000000000000000000000000000000000000111111110000,
		56'b00000000000000000000000000000000000000000000111111110000,
		56'b00000000000000000000000000000000000000000000111111110000,
		56'b00000000000000000000000000000000000000000000011111110000,
		56'b00000000000000000000000000000000000000000000000010000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 5
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000001111111111000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111111110000000000000000000000,
		56'b00000000000000000000000011111111111111110000000000000000,
		56'b00000000000000000000000011111111111111111111000000000000,
		56'b00000000000000000000000011111111111111111111000000000000,
		56'b00000000000000000000000001111111111111111111000000000000,
		56'b00000000000000000000000001111110011111111111000000000000,
		56'b00000000000000000000000001111110000000000110000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111110000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111110000000000000000000000,
		56'b00000000000000000000000001111111111000000000000000000000,
		56'b00000000000000000000000001111111111100000000000000000000,
		56'b00000000000000000000000000111111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111100011111110000000000000000,
		56'b00000000111111000000000000111110011111110000000000000000,
		56'b00000001111111111000000000111110001111111000000000000000,
		56'b00000001111111111110000000111110000111111100000000000000,
		56'b00000001111111111111110000111110000001111110000000000000,
		56'b00000000111111111111111100111110000001111110000000000000,
		56'b00000000000000111111111111111110000000111111000000000000,
		56'b00000000000000001111111111111110000000011111000000000000,
		56'b00000000000000000011111111111110000000011111000000000000,
		56'b00000000000000000000011111111110000000011111100000000000,
		56'b00000000000000000000000011111110000000001111100000000000,
		56'b00000000000000000000000000111100000000001111100000000000,
		56'b00000000000000000000000000000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000111110000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000011111000000000,
		56'b00000000000000000000000000000000000000000011111100000000,
		56'b00000000000000000000000000000000000000000001111111100000,
		56'b00000000000000000000000000000000000000000001111111110000,
		56'b00000000000000000000000000000000000000000001111111110000,
		56'b00000000000000000000000000000000000000000000111111100000,
		56'b00000000000000000000000000000000000000000000011111000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 6
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111100000000000000000000,
		56'b00000000000000000000000000001111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000011111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000011111111111100000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000001111111111000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000000111111000000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111000000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000000111111111000000000000000000000,
		56'b00000000000000000000000000111111111100000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000000111111111111110000000000000000,
		56'b00000000000000000000000001111111111111111000000000000000,
		56'b00000000000000000000000001111101111111111000000000000000,
		56'b00000000000000000000000001111111111111111000000000000000,
		56'b00000000000000000000000001111111111110000000000000000000,
		56'b00000000000000000000000000111111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111110000000000000000000,
		56'b00000000000000000000000000011111111100000000000000000000,
		56'b00000000000000000000000000011111111100000000000000000000,
		56'b00000000000111111110000000011111111110000000000000000000,
		56'b00000000000111111111100000011111111110000000000000000000,
		56'b00000000000111111111111000001111111111000000000000000000,
		56'b00000000000111111111111110001111111111100000000000000000,
		56'b00000000000011111111111111101111111111110000000000000000,
		56'b00000000000000000011111111111111101111110000000000000000,
		56'b00000000000000000000111111111111110111111000000000000000,
		56'b00000000000000000000001111111111110011111000000000000000,
		56'b00000000000000000000000011111111110011111000000000000000,
		56'b00000000000000000000000000111111110011111000000000000000,
		56'b00000000000000000000000000001111110001111100000000000000,
		56'b00000000000000000000000000000001100001111100000000000000,
		56'b00000000000000000000000000000000000001111100000000000000,
		56'b00000000000000000000000000000000000001111110000000000000,
		56'b00000000000000000000000000000000000000111110000000000000,
		56'b00000000000000000000000000000000000000111110000000000000,
		56'b00000000000000000000000000000000000000111111000000000000,
		56'b00000000000000000000000000000000000000011111000000000000,
		56'b00000000000000000000000000000000000000011111000000000000,
		56'b00000000000000000000000000000000000000011111000000000000,
		56'b00000000000000000000000000000000000000001111100000000000,
		56'b00000000000000000000000000000000000000001111111100000000,
		56'b00000000000000000000000000000000000000001111111100000000,
		56'b00000000000000000000000000000000000000000111111100000000,
		56'b00000000000000000000000000000000000000000111111100000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,

		//Page 7
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111000000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000111111111000000000000000000000000,
		56'b00000000000000000000000111111111110000000000000000000000,
		56'b00000000000000000000000111111111111100000000000000000000,
		56'b00000000000000000000000111111111111111100000000000000000,
		56'b00000000000000000000000111111111111111111000000000000000,
		56'b00000000000000000000000111111111111111111111000000000000,
		56'b00000000000000000000000111111110011111111111100000000000,
		56'b00000000000000000000000011111110000011111111100000000000,
		56'b00000000000000000000000011111110000000111111100000000000,
		56'b00000000000000000000000011111100000000000111000000000000,
		56'b00000000000000000000000011111100000000000000000000000000,
		56'b00000000000000000000000011111110000000000000000000000000,
		56'b00000000000000000000000011111110000000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000011111111000000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000000111111110000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000001100000011111111100000000000000000000,
		56'b00000000000000000111111111011111111100000000000000000000,
		56'b00000000000000001111111111111111111110000000000000000000,
		56'b00000000000000011111111111111111111111000000000000000000,
		56'b00000000000000011111111111111111111111000000000000000000,
		56'b00000000000000011111001111111111111111100000000000000000,
		56'b00000000000000011110000000111111111111100000000000000000,
		56'b00000000000000000000000000000111111111100000000000000000,
		56'b00000000000000000000000000000111110110000000000000000000,
		56'b00000000000000000000000000000111110000000000000000000000,
		56'b00000000000000000000000000000111110000000000000000000000,
		56'b00000000000000000000000000000111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000001111000000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000011111000000000000000000000000,
		56'b00000000000000000000000000011111110000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000011111111000000000000000000000,
		56'b00000000000000000000000000001111110000000000000000000000,

		//Page 8
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000111111000000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000001111111111111000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000001111111000000000000000000000,
		56'b00000000000000000000000000001111100000000000000000000000,
		56'b00000000000000000000000000011111100000000000000000000000,
		56'b00000000000000000000000000111111100000000000000000000000,
		56'b00000000000000000000000001111111100000000000000000000000,
		56'b00000000000000000000000011111111100000000000000000000000,
		56'b00000000000000000000000111111111100000000000000000000000,
		56'b00000000000000000000000111111111100000000000000000000000,
		56'b00000000000000000000001111111111100000000000000000000000,
		56'b00000000000000000000011111111111100000000000000000000000,
		56'b00000000000000000000111111011111100000000111110000000000,
		56'b00000000000000000000111111011111100001111111111000000000,
		56'b00000000000000000001111110011111111111111111111000000000,
		56'b00000000000000000001111100011111111111111111110000000000,
		56'b00000000000000000001111100111111111111111111100000000000,
		56'b00000000000000000011111000111111111111111000000000000000,
		56'b00000000000000000011111000111111111110000000000000000000,
		56'b00000000000000000011111000111111100000000000000000000000,
		56'b00000000000000000011111000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110000111110000000000000000000000000,
		56'b00000000000000000111110001111110000000000000000000000000,
		56'b00000000000000000111110001111100000000000000000000000000,
		56'b00000000000000001111100001111110000000000000000000000000,
		56'b00000000000000001111100001111111000000000000000000000000,
		56'b00000000000000001111100001111111110000000000000000000000,
		56'b00000000000000001111100001111111111000000000000000000000,
		56'b00000000000000001111000001111111111110000000000000000000,
		56'b00000000000000000000000001111111111111000000000000000000,
		56'b00000000000000000000000001111101111111110000000000000000,
		56'b00000000000000000000000000111100111111111000000000000000,
		56'b00000000000000000000000001111100001111111110000000000000,
		56'b00000000000000000000000000111110000011111111000000000000,
		56'b00000000000000000000000000111111111111111111000000000000,
		56'b00000000000000000000000000111111111111111111000000000000,
		56'b00000000000000000000000011111111111111111111000000000000,
		56'b00000000000000000000000111111111111111111100000000000000,
		56'b00000000000000000000000111111111111110000000000000000000,
		56'b00000000000000000000001111111111000000000000000000000000,
		56'b00000000000000000000001111111110000000000000000000000000,
		56'b00000000000000000000001111111110000000000000000000000000,
		56'b00000000000000000000000111111110000000000000000000000000,
		56'b00000000000000000000000011111110000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000001111100000000000000000000000000,
		56'b00000000000000000000000011111000000000000000000000000000,
		56'b00000000000000000000000011111000000000000000000000000000,
		56'b00000000000000000000000111110000000000000000000000000000,
		56'b00000000000000000000000111110000000000000000000000000000,
		56'b00000000000000000000000111110000000000000000000000000000,
		56'b00000000000000000000001111100000000000000000000000000000,
		56'b00000000000000000000001111100000000000000000000000000000,
		56'b00000000000000000000001111100000000000000000000000000000,
		56'b00000000000000000000011111000000000000000000000000000000,
		56'b00000000000000000000011111000000000000000000000000000000,
		56'b00000000000000000000111111100000000000000000000000000000,
		56'b00000000000000000000111111110000000000000000000000000000,
		56'b00000000000000000000111111110000000000000000000000000000,
		56'b00000000000000000000111111110000000000000000000000000000,
		56'b00000000000000000000000111000000000000000000000000000000,

		//Page 9
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000,
		56'b00000000000000000000000000001111111100000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111000000000000000000,
		56'b00000000000000000000000000111111111111000000000000000000,
		56'b00000000000000000000000000011111111111000000000000000000,
		56'b00000000000000000000000000011111111110000000000000000000,
		56'b00000000000000000000000000001111111000000000000000000000,
		56'b00000000000000000000000000111111100000000000011000000000,
		56'b00000000000000000000000001111111100000000000111100000000,
		56'b00000000000000000000000111111111110000000001111110000000,
		56'b00000000000000000000011111111111110000000011111100000000,
		56'b00000000000000000001111111111111111000000111111100000000,
		56'b00000000000000000111111111111111111000001111111000000000,
		56'b00000000000000001111111110011111111100011111110000000000,
		56'b00000000000000001111111100011111111100111111100000000000,
		56'b00000000000000001111110000011111111111111111000000000000,
		56'b00000000000000001111100000011111111111111110000000000000,
		56'b00000000000000001111100000011111011111111100000000000000,
		56'b00000000000000001111100000011111011111111000000000000000,
		56'b00000000000000001111100000011110001111110000000000000000,
		56'b00000000000000001111000000111110001111100000000000000000,
		56'b00000000000000001111000000111110000111000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000000111110000000000000000000000000,
		56'b00000000000000011111000001111100000000000000000000000000,
		56'b00000000000000011111000001111100000000000000000000000000,
		56'b00000000000000011110000001111111100000000000000000000000,
		56'b00000000000000001100000001111111111100000000000000000000,
		56'b00000000000000000000000001111111111111100000000000000000,
		56'b00000000000000000000000001111111111111111100000000000000,
		56'b00000000000000000000000001111111111111111111100000000000,
		56'b00000000000000000000000001111100011111111111110000000000,
		56'b00000000000000000000000001111100000011111111110000000000,
		56'b00000000000000000000000001111100000000111111110000000000,
		56'b00000000000000000000000001111000000000111111110000000000,
		56'b00000000000000000000000011111000000001111111000000000000,
		56'b00000000000000000000000011111000000111111110000000000000,
		56'b00000000000000000000000011111000001111111100000000000000,
		56'b00000000000000000000000011111000011111111000000000000000,
		56'b00000000000000000000000011111000111111100000000000000000,
		56'b00000000000000000000000011111011111111000000000000000000,
		56'b00000000000000000000000011111111111110000000000000000000,
		56'b00000000000000000000000011111111111100000000000000000000,
		56'b00000000000000000000000111111111110000000000000000000000,
		56'b00000000000000000000000111111111111000000000000000000000,
		56'b00000000000000000000001111110111111000000000000000000000,
		56'b00000000000000000000011111100011111000000000000000000000,
		56'b00000000000000000000111111000001110000000000000000000000,
		56'b00000000000000000000111111000000000000000000000000000000,
		56'b00000000000000000001111110000000000000000000000000000000,
		56'b00000000000000000011111100000000000000000000000000000000,
		56'b00000000000000000111111000000000000000000000000000000000,
		56'b00000000000000001111111000000000000000000000000000000000,
		56'b00000000000000011111110000000000000000000000000000000000,
		56'b00000000000000011111100000000000000000000000000000000000,
		56'b00000000000000111111000000000000000000000000000000000000,
		56'b00000000000001111110000000000000000000000000000000000000,
		56'b00000000000001111110000000000000000000000000000000000000,
		56'b00000000000001111110000000000000000000000000000000000000,
		56'b00000000000001111111000000000000000000000000000000000000,
		56'b00000000000000111111000000000000000000000000000000000000,
		56'b00000000000000011111000000000000000000000000000000000000,
		56'b00000000000000001110000000000000000000000000000000000000,
		56'b00000000000000000000000000000000000000000000000000000000

        };

	assign data = ROM[addr];

endmodule  


module cover_rom ( input [9:0] addr, output [639:0] data);

	//parameter ADDR_WIDTH = 9;
	parameter ROM_LENGTH = 480;	//
	parameter DATA_WIDTH = 640;
				
	// ROM definition:
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {
		
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000001111110000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000111111100000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000001111111000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000111111100000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011111111000000000000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000111111111000000000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000001111111100000000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000011111110000000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000111111100000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000011111110000000111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000001111111100000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000011111111000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000001111111100111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011111110111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000111111111100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000011111111100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000001111111100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000011111110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000001111110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000111111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000011111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000011111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000010000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111111100000000000011111111111111111110000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000001111111111111111111111100000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011110000000000001111111111111111111111100000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000001111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000001111000000000000001111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000001111000000000000001111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000001111000000000000001111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111000000000000001111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111000000000000001111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111000000000000000111100000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111111000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111100000000000000111100000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000011111000000011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000000000111100000000000000000000000000000000000011000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000111100000111111100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000001111000000000001111100000000000000111100000000000000000000000011111111111111100000000000001110000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000111000000000111100011111110000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000001111000000000001111111111111111111111100000000000000000000000011111111111111100000000000001110000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000001111000000000011111111111000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000001111000000000001111111111111111111111110000000000000000000000111111111111111100000000000001110000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000001111000000000001111111110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000001110111111111110000000000000000000000000000000000000000000111000000000001111111111111111111111110000000000000000000000111111000000111100000000000001110000000000000000000000000000000000000000000000000000000000011111111000001111111111000000000000000000000000000000000000000000000000000000000001110000000000001111111000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000001110001111111111000000000000000000000000000000000000000000111000000000000111111111111111111111110000000000000000000000011110000000011100000000000001110000000000000000000000000000000000000000000000000000000000111111000000000011111111110000000000000000000000000000000000000000000000000000000001110000000000001111110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000001110000000111111000000000000000000000000000000000000000000111000000000000001000000001111111111100000000000000000000000011110000000011100000000000001110000000000000000000000000000000000000000000000000000000000111100000000000000111111111000000000000000000000000000000000000000000000111111111001110000000000000111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000001110000000011111000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000011110000000011100000000000001110000000000000000000000000000000000000000000000000000000001111000000000000000000111111000000000000000000000000000000000000000001111111111111111110000000000000111100000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000011100000000111111000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000011110000000111100000000000001110000000000000000000000000000000000000000000001111100000011110000000000000000000001111100000000000000000000000000000000000000111111111111111111100000000000000111110000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000011100000000111111000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000011110000000111100000000000001110000000000000000000000000000000000000000001111111111000111100000000000000001110000111110000000000000000000000000000000000001111111110000001111100000000000001111111000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000011100000000111111100000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000011110000000011100000000000001110000000000000000000000000000000000000000011111111111111111100000000000000111111100111110000000000000000000000000000000000011111110000000000011110000000000011111111110000000000000000000111000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000111111000000001111110000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000011110000000011110000000000001110000000000000000000000000000000000000001111111111111111111100000000000000111111110011111000000000000000000000000000000000111111000000000000001111000000000111111111111100000000000000000111000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000011111111000000000000000000000000000000000111000000000000000000000000000000111111000000000111111100000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000011110000000011110000000000001110000000000000000000000000000000000000011111000000011111111000000000000000111111110011111000000000000000000000000000000001111100000000000000001110000000001111000001111100000000000000001111000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001111111110000000000000000000000000000011111111100000000000000000000000000111111000000000011111111000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000011111000000011110000000000001110000000000000000000000000000000000000011110000000000111110000000000000000111101111001111000000000000000000000000000000001111000000000000000000000000000001111000000011110000000000000001111000000000000000000000000000000000000000000000000000111100111111000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000111111111000000000000000000000000000011111111110000000000000000000000000111110000000000000111111100000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000001111000000011111000000000001111000000000000000000000000000000000000111110000000000000000000000000000001111101111001111000000000000000000000000000000011110000000000000000000000000000011110000000001110000000000000001110000000000000000000000000000000000000000000000000000111000011111000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000001111111111000000000000000000000000011111111111111111000000000000000000011110000000000000011111111000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000001111000000011111000000000001111000000000000000000000000000000000000111100000000000000000000000000000001111000111001111100000000000000000000000000000011110000000000000000000000000000011100000000001110000000000000001110000000000000000000000000000000000000000000000000001111000001111110000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000011111111110000000000000000000000011100011111111111100000000000000000011100000000000000000111111111000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000001111000000001111000000000001111000000000000000000000000000000000001111100000000000000000000000000000001111000111000111100000000000000000000000000000111100000000000000000000000000000001000000000001110000000000000011110000000000000000000000000000000000000000000000000011110000000111111100000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000111111111110000000000000000000011100000011111111100000000000000000111100000000000000000111111111100000000000000000000000000000011110000000000000000000000000000000000000000000000000000000001111000000001111000000000001111000000000000000000000000000000000001111000000000000000000000000000000001111111111000111100000000000000000000000000000111100000000000000000000000000000000000000000011100000000000000111100000000000000000000000000000000000000000000000000111100000000001111110000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000111111111100000000000000000011100000000111111100000000000000000111100000000000000011111111111100000000000000000000000000000011110000000000000000000000000000000000000000000000000000000001111100000001111000000000001111000000000000000000000000000000000001111000000000000000000000000000000001111111111000111100000000000000000000000000000111100000000000000000000000000000000000000000011100000000000000111100000000000000000000000000000000000000000000000001111000000000000011111000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001111111110000000000000000011100000001111111000000000000000000111000000000000000111111111111000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000001111100000001111000000000001111000000000000000000000000000000000001111000000000000000000000000000000001111111111000111100000000000000000000000000000111100000000000000000000000000000000000000000011100000000000001111000000000000000000000000000000000000000000000000011110000000000000001111100000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000011111111100000000000000111100000001111111100000000000000001111000000000000111111111111110000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000111100000001111000000000001111000000000000000000000000000000000001111100000000000000000000000000000000111111110000111100000000000000000000000000000011110000000000000000000000000000000000000000000000111000000011110000000000000000000000000000000000000000000000000111100000000000000000111110000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111100000000000000000000000000000000000111111111000000000000111100000000111111111000000000000001111011111110000111111110000000000000000000000000000000000000001110000000000000000000000000000000000001111111111111111111111111111111111111111111111011111000000000000000000000000000000000000111100000000000000000000000000000000000011100000111100000000000000000000000000000011110000000000000000000000000000000000000000000001111000011111110000000000000000000000000000000000000000000000001111000000000000000000011111000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111100000000000000000000000000000000000001111111100000000000111111000000001111111110000000000001111111111111001111110000000000000000000000000000000000000000001111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111000000000000000000000000000000000000000000111100000000000000000000000000000001111000000000000000000000000000000000000000000000111100011111100000000000000000000000000000000000000000000000001111000001111000000000001111110000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000111111110000000000111111100000000011111111100000000001111111111111000111100000000000000000000000000000000000000000001111000000000000000000011111111111111111100000000000000000000000000000000111000000011111111111111111100000000000000000000000000011111111111100000000000000000000000000000000000011111100000000000000000000000000001111000000001000000000000000000000000000000000000111110011111100000000000000000000000000000000000000000000000011110000011111000000000000111111000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000011111111100000000000111111100000000000111111110000000001111110001111100111100000000000000000000000000000000000000000001111000000000011111111111100000000000000000000000000000000000000000000000000000000000000110000000011111111111100000000000000000001111111111111000000000000000000000000000000000011111110000000000000000000000000000111100001111110000000000000000000000000000000000011111000111110000000000000000000000000000000000000000000000111100000111111100000000000001111100000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000001111111111000000000000111111100000000000001111111110000001111100000111100011100000000000000000000000000000000000000000001111001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000011111111111111111100000000000000000000000000001111111100000000011110000000000000011100111111111100000000000000000000000000000000001111000001111000000000000000000000000000000000000000000001111000001111111111000000000000111110000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000111111111000000000000001111111100000000000000011111111000000111000000111100011110000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000001111111111111111000000000000000000000000011111111000001111110000000000000000001111111111000000000000000000000000000000000001111000000111100000000000000000000000000000000000000000011110000001110011111100000000000011111000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110111100000000000000000000000000000011111111000000000000000001111111100000000000000001111111000000000000000011110011110000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000111111111111111111100000000000000000000000111111110011111110000000000000000001111100000000000000000000000000000000000000000111100000111100000000000000000000000000000000000000000111100000011110000111100000000000001111100000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000111100000000000000000000000000000111111100000000000000000001110011100000000000000001111111000000000000000011110001111000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000111111111111111111111110000000000000000000001111110011111100000000000000000001111000000000000000000000000000000000000000000111100000011100000000000000000000000000000000000000001111000000111100000111110000000000000111110000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000011111111000000000000000000000000011100000000000000011111110000000000000000001111001111000000000000000000000000000111111110000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000111111111111100000000000000000000011111000110000000000000000000011110000000000000000000000000000000000000000000111100000011100000000000000000000000000000000000000011110000001111000000111100000000000000011111000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000011111100000000000000000000000000011100000000000011111111100000000000000000001111001111100000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000011111111111111000000000000000001111000000000000000000000000011110000000000000000000000000000000000000000001111000000011100000000000000000000000000000000000000111110000011110000001111100000000000000001111100000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000111111000000000000000000000000000011100000000000111111110000000000000000000000111000111100000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000001111111111110000000000000001111000000000000000000000000011110000000000000000000000000000000000000000111111000000011100000000000000000000000000000000000001111100000011110000011111000000000000000000111110000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000001111110000000000000000000000000000011100000110000111111100000000000000000000000111100111110000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000111111111110000000000001111000111000000000000000000011110000000000000000000000000000000000011111111110000000011100000000000000000000000000000000000001111000000011100000111110000000000000000000011111100000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000001111000000000000000000000000000000011100001111000111110000000000000000000000000111110011110000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000011111111000000000001111001111100000000000000000011110000000000000000000000000000000000011111111000000000011100000000000000000000000000000000000011110000000011110000111100000000000000000000000111100000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000001111000000000000000000000000000000011100111111100011111000000000000000000000000011110011111000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000001111111111100000011111000111110000000000000000001110000000000000000000000000000000000011111110000000000111100000000000000000000000000000000000111100000000011111001111000000000000000000000000011110000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000111100000000000000000000000000000011101111111100011111000000000000000000000000011110001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111111100011110000111100000000000000000001110000000000000000000000000000000000011111100000000000111100000000000000000000000000000000001111100000000001111111110000000000000111100000000001111000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000011000000111110000000000000000000000000000011111111111110001111100000000000000000000000001111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111111111110011000000000000000000000001111000000000000000000000000000000000000000000000000001111000000000000000000000000000000000011111000000000000111111110000000000001111110000000000111110000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000011110111100000011111000000000000000000000000000011111110011110001111100000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000111111111111100111100000000000000000000001111100000000000000011000000000000000000000000000000001111000000000000000000000000000000000111110000000000000011111110000000000011111111000000000011111000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111111111110000011111000000000000000000000000000011111100001111000111110000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100001111111111111100111100000000000000000000000111100000000000000111000000000000000000000000000000011110000000000000000000000000000000000111100000000000000000110000000000000111111111100000000001111000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000011111110011110000001111100000000000000000000000000111111000001111100011110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000011100000000000000000000000111111000000000000111000000000000000000000000000000111100000000000000000000000000000000001111000000000000000000000000000000001111100111100000000000111100,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000111111000011111000000111100000000000000000000000000011110000001111100011111000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000011100000000000000000000000011111100000000001111000000000000000000000011111111111100000000000000000000000000000000011111000001111110000000000000000000001111000011110000000000011110,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011111110000001111000000111110000000000000000000000000011100000000111110001111100000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001100000000000000000000000001111111111000011110000000000000000000000011111111110000000000000000000000000000000000111110000001111110000000000000000000011110000011110000000000011111,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000111111100000000111100000011111000000000000000000000000000000000000111110001111100000000000011111100000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000011111111000011110000010000000000000000011111111100000000000000000000000000000000001111100000011111111000000000000000000111100000011110000000000001111,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001111110000000000111100000011111000000000000000000000000000000000000011111000111110000000001111000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000111111000111100000111000000000000000001111000000000000000000000000000000000000011111000000011110111100000000000000001111000000011110000000000001111,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011111100000000000011111000001111100000000000000000000000000000000000001111000011111000011111110000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000111100001110000000000000000001111000000000000000000000000000000000000011110000000111100111111000000000000001111000000111100000000000001111,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001111111000000000000011111000001111110000000000000000000000000000000000001111100011111101111110000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111000011110000000000000000001111000000000000000000000000000000000000111100000000111000011111000000000000011110000001111100000000000011111,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111110000000000000001111100000111110000000000000000000000000000000000000111100001111111110000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000011111000011100000000000000000001111000000000000000000000000000000000001111100000001110000001111000000000000011110000011111000000000000011110,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000111100000011111000000000000000000000000000000000000111110001111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011110000111100000000000000000001111000000000000000000000000000000000011111000000011110000011110000000000000011110000111110000000000000111100,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111110000001111000000000000000000000000000000000000011111011111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000111100001111000000000000000000001111000000000000000000000000000000000011110000000111100000111100000000000000011111001111000000000000001111000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000011110000001111100000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000001111100001111000000000000000000001111000000000000000000000000000000000111100000001111000001111000000000000000001111111111000000000000011110000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000011111000000111110000000000000000000000000000000000011111110000000000000000000000000000000000000000000000100000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000001111000011110000000000000000000001111000000000000000000000000000000001111000000011111000011110000000000000000000111111110000000000000111110000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000001111000000111111000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000011111000111110000111000000000000011110000000000000000000000000000000011111000000011110000111100000000000000000000001111100000000000001111100000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011111100000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011110000111100000111100000000001111100000000000000000000000000000000111110000000001111111111000000000000000000000000110000000000000011111000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000001111100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000111110001111000000111110000000011111000000000000000000000000000000000111100000000000111111111000000000001110000000000000000000000000011110000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000111110000000000000000000000001111110000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000111100001111000000011111111111111111000000000000000000000000000000001111000000000000011111110000000000011111110000000000000000000000111100000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000001111000011110000000011111111111111100000000000000000000000000000000011111000000000000000111100000000000111111111000000000000000000001111100000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011111000000000000000000011111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000011111000111100000000001111111111110000000000000000000000000000000000111110000000000000000000000000000001111001111100000000000000000011111000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000001111100000000000000001111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000011110000111100000000000001111110000000000000000000000000000000000000111100000011100000000000000000000011110000111110000000000000000111110000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000111110000000000000111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000011110000111100001111000000000000000000000000000000000000000000000000000000001111000000111110000000000000000000111100000011110000000000000001111100000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000111110000000000011111000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000001111100111100001111000000000000000000000000000000000000000000000000000000011111000001111111100000000000000001111000000011110000000000000011111000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000011111000000001111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000011111111000011110000000000000000000000000000000000000000000000000000000111110000011111111110000000000000011111000000111100000000000000111110000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011111100000111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000111111000011100000000000000000000000000000000000000000000000000000001111100000111110011110000000000000111110000001111100000000000001111100000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000001111100001111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000001111000111100000000000000000000000000000000000000000000000000000001111000001111100001110000000000000111100000001111000000000000011111000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000111110111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000011110000001111000011110000000000000111110000011110000000000000011110000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000011111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000111110000011110000011110000000000000011111100011100000000000000111100000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000011111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000001111100000111110000111100000000000000001111111111100000000000001111100000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000001111000000111100001111100000000000000000011111111000000000000011111000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110001111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011101111000000000000000000000000000000000000000000000000011110000001111000001111000000000000000000000111110000000000000111110000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000111100000011110000011110000000000111100000000011110000000000001111100000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111100000011110000111100000000001111110000000001100000000000011111000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000011111000000011111111111000000000011111111000000000000000000000011110000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000111110000000001111111111000000000111111111000000000000000000000111110000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111110000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000111100000000000001111110000000000111100111100000000000000000001111100000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111110000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000001111000000000000000111000000000001111000111111000000000000000011111000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110001111111111110000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000011110000000011100000000000000000011110000011111000000000000000111110000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001111111000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100011111111111110000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000111110000001111110000000000000000111110000001111000000000000001111100000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111100000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000011111111111110000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000001111100000011111111000000000000001111100000001111000000000000011111000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000011111111111110000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111000000111101111000000000000001111000000011110000000000000011110000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011111000001111100111100000000000011110000000111100000000000000111100000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110011110000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000111110000011111000111100000000000111111000001111000000000000001111100000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110111111000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000001111100000011110000111100000000000111111100011110000000000000011111000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000011111111110001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011111000000111100000111000000000000001111110111100000000000000111110000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000011111000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000011110000001111000001111000000000000000011111111000000000000000111100000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000011111000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000001111110000001111000011110000000000000000001111111000000000000001111100000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000001111111110000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001111100000011111000111110000000001110000000111110000000000000011111000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000011111111110000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011111000000011111101111000000000011111000000011110000000000000111110000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000111110011110000000000000000000000000001100011111111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000111110000000001111111110000000000111111100000000000000000000001111100000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000001111100001111000000000000000000000000011110011111110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000011111100000000000000000000001100000000000000000000000000000111111111110000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111100000000000011111100000000001111111100000000000000000000011111000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000011111000001111100000000000000000000000011111111111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000000111111100000000000000000000011111000000000000000000000000000000111111111000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000001111100000000011110111110000000000000000000111111000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000001111110000000111110000000000000000000000111111111111110000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000111111100000000000000000000111111000000000000000011111111111110011111111100000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000111100011111100000000000000001111110000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000011111100000000011111000000000000000000000111111111111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000111111100000000000000000000111111000000000000001111111111111111101111111110000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000001111000001111110000000000000001111100000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000111111000000000001111000000000000000000000011111111011111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111011111111111111111111110000000000000000001111111100000000000000000000111111000000000000011111111111111111110111111111000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000011110000000111100000000000000011111000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000111100000000000000111100000000000000000000011110000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111100000000000000000001111111100000000000000000000111111000000000000111111111111111111111011111111000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101110000000000000000000000011100000000111100000000000000111110000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000011111000001110000000011110000000000000011110011110000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000111111111111111111100000000000000000001111111100000000000000000000111111000000000001111111111111111111111111111111100000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111000000000000000000000111100000001111100000000000001111100000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000111111000011111000000011111000000000000011111111110000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111000000000000000000001111111100000000000000000000111111000000000001111111111111111111111111111111110000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000111110000011111000000000000011111100000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000111110000111111100000001111100000000000011111111110000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111011111111111111111110000000000000000000001111111100000000000000000000111111100000000011111111111111111111111111111111110000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000111111100111110000000000000011111000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000001111100001111111100000000111110000000000001111111100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000001111111110000000000000000000111111100000000011111111111111111111111111011111110000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000001111111111100000000000000111110000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000011111000011111111100000000011111000000000000111110000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000001111111110000000000000000001111111100000000111111111111111111111111111111111110000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000111111111000000000000000111100000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000011110000111111011110000000001111100000000000111111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000001111111110000000000000000001111111100000000111111111110000001111111111101111110000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000001111110000000000000001111000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000111100000111110011110000000000111100000000000011111100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000001111111110000000000000000001111111100000000111111111100000000011111111100111110000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111110000000000000011111000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000001111100000111111111100000000000111110000000000001111101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000001111111110000000000000000001111111100000000111111111000000000001111111110011100000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000011100000000000000111110000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000011111000000011111111000000000000011111000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000001111111110000000000000000001111111100000001111111111000000000001111111110000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000001111100000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000111110000000001111110000000000000001111100000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111110000000000000001111111110000000000000000001111111100000001111111110000000000000111111111000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000011111000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000001111100000000000111100000000000000000111110000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111100000000000001111111110000000000000000001111111100000001111111110000000000000111111111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000011110000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000011111000000000000001000000000000000000011111100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100001111111111111111110000000000001111111110000000000000000001111111100000011111111100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000111110001111100000000000000000000000000001111110000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000111111111111111111000000000000111111110000000000000000001111111100000011111111100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000001111100000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000001111100011111100000000000000000000000000001111110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000011111111111111111100000000000111111111000000000000000001111111100000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000001111000111111110000000000000000000000000011111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000011111111111111111110000000000111111111000000000000000011111111100000011111111000000000000000011111111100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000011110000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000011111001111111110000000000000000000000000111111110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000001111111111111111111000000000111111111100000000000000011111111100000011111111000000000000000011111111100000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000111110000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000111100001111101111100000000000000000000001111110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000111111111111111111100000000111111111110000000000000011111111000000011111111000000000000000001111111100000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000001111100000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000001111100011111000111100000000000000000000011111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000111111111111111111110000000011111111110000000000000011111111000000111111111000000000000000001111111100000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000011111000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000011110000011111001111100000000000000000000111111000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000011111111111111111111000000011111111111000000000000111111111000000111111110000000000000000000111111100000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011110000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000111110000011111011111100000000000000000000111111100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000001111111111111111111100000011111111111100000000001111111111000000111111110000000000000000000111111100000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000111100000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000001111100000011111111111000000000000000000011111111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000001111111111111111111110000011111111111110000000001111111111000000111111110000000000000000000111111100000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111100000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000011111000000001111111110000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000111111111111111111110000011111111111111000000111111111111000000111111110000000000000000000111111100000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000011111000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000111110000000000111111100000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000011111111111111111111000001111111111111111111111111111111000000111111110000000000000000000111111100000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111110000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000001111100000000000011111000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000001111111111111111111100001111111111111111111111111111110000000111111110000000000000000000111111100000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000111100000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000011111000100000000001110000000000000000000111111011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000001111111111111111111110001111111111111111111111111111110000000111111110000000000000000000111111100000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111100000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000111110011111000000000000000000000000000001111110001111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111110000000000000000000111111111111111111111000111111111111111111111111111110000000111111110000000000000000000111111100000000000000000011111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001110011111000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000001111100111111100000000000000000000000000011111100001110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111110000000000000000000111111111111111111111000111111111111111111111111111100000000111111100000000000000000000111111100000000000000000011111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000011111000111111110000000000000000000000000111111000011100000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111000000000000000000011111111111111111111100011111111111111111111111111100000000111111100000000000000000000111111100000000000000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000111110001111111111000000000000000000000001111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000001111111111111111111000001111111111111111111111111000000000111111100000000000000000000111111100000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000001111100001111001111100000000000000000000011111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000001111111111111111111000000111111111111111111111110000000000111111000000000000000000000111111100000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000011111000011111000111100000000000000000000111111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000111111111111111110000000011111111111111111111100000000000011110000000000000000000000011111000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000111110000011111001111100000000000000000001111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000011111111111111100000000000111111111111111111000000000000000000000000000000000000000001110000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000111100000011111111111100000000000000000011111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000001111111111111000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000001111000000001111111111000000000000000000011111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000111111111110000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000011111000000000111111110000000000000000001111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000111110000000000011111100000000000000000011111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000001111000000000000000000000000000000000000000000,
		640'b00000000000000000000000000001111100000000000000111000000000000000000011111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000011111000000000000000000000000000000000000000000,
		640'b00000000000000000000000000011111000000000000000000000000000000000000111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111000000000000000000000000000000000000000000,
		640'b00000000000000000000000000111110000111100000000000000000000000000001111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000111111100000011000000000000000000000000000000000,
		640'b00000000000000000000000000111100000111110000000000000000000000000011111000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111111100111111100000000000000000000000000000000,
		640'b00000000000000000000000001111100001111111100000000000000000000000111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011111111111111111100000000000000000000000000000000,
		640'b00000000000000000000000011111000011111111110000000000000000000001111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000,
		640'b00000000000000000000000111100000011110111110000000000000000000011111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111111111100000000000000000000000000000000,
		640'b00000000000000000000000111100000111100011110000000000000000000011111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100001111001111000000000000000000000000000000000,
		640'b00000000000000000000001111000000111110111100000000000000000000111110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001000000000000000100000000000000000110000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000001111000000000000000000000000000000000,
		640'b00000000000000000000001111000000011111111100000000000000000001111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011111110000000001110000000000000011111000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011111000000000000000000000000000000000,
		640'b00000000000000000000000111100000001111111000000000000000000011111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000001000000001100000000000111110000011111111000000001110000000000001111111000011111100000000000000000000000000111100000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000011111000001100000000000000000000000000,
		640'b00000000000000000000000111110000000011110000000000000000000111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000001111111000001111111000001111100000111100000000001111000000011100111100000011111000000000111110000000011000000000000111111111111000011111111000000000000011110111111111111100000110000000011111111001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111000011110000000000000000000000000,
		640'b00000000000000000000000011111100000001110000000000000000001111110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110001111111100001111111000011111000001111100000000001100000000011100011100000011111100000001111000000000011000000000000111111111111001111111111100000000001111110111111111111100001111000000011111111101111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000011111111111110000000000000000000000000,
		640'b00000000000000000000000001111110000000000000000000000000001111100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001110001110011110001110000000111100000011100000000000011110000000011100011100000111011100000001110000000000011000000000000000001110000001110000001110000000001110000000001110000000001111000000001100011100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000001111111111110000000000000000000000000,
		640'b00000000000000000000000000111111000000000000000000000000011111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000110001110001110001110000000111000000011100000000000001111000000011100011100000111001110000011100000000000011000000000000000001110000011100000001110000000011110000000001110000000011111100000001100011100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111111111110000000000000000000000000,
		640'b00000000000000000000000000011111110000000000000000000000111110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001110001110011100001110000000111100000011110000000000001111110000011100111000001110001110000011100000000000011111100000000000001110000011100000000111000000001111000000001110000000011001110000001100011100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111111100000000000000000000000000,
		640'b00000000000000000000000000000111111000000000000000000001111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001110001110111100001111111000011111000011111000000000000011111000011101111000001110111111000011100000000000011111100000000000001110000011000000000111000000001111100000001110000000111001110000001100111000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000111111111100000000000000000000000000,
		640'b00000000000000000000000000000111111100000000000000000011111100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100001111111000001111111000001111100000111110000000000000111000011111110000011111111111000011100000000000011000000000000000001110000111000000000111000000000011110000001110000000111111111000001101110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111110111100001111100000000000000000,
		640'b00000000000000000000000000000001111110000000000000000111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000001110111000001110000000000011100000001110000000000000111000011111000000011111111111100011100000000000011000000000000000001110000111000000000110000000000001111000001110000001111111111000001101111000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011111100111111111111100000000000000000,
		640'b00000000000000000000000000000000111111000000000000001111110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000001110011100001110000000000001100000001110000000000000111000011100000000111000000011100011110000000000011000000000000000001110000011100000001110000000000000111000001110000001111111111100001100111100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011111000011111111111100000000000000000,
		640'b00000000000000000000000000000000011111100000000000011111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001110001110001110000000000011100000011110000000000001111000011100000000111000000001110001111000000000011000000000000000001110000011110000011100000000000001110000001110000011100000011110001100011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000011111111111100000000000000000,
		640'b00000000000000000000000000000000001111110000000000111111110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001110001111001111111000011111000001111100000000001111110000011100000001110000000001111000111111111100011111110000000000001110000001111111111100000000001111110000001110000111000000001110001100001111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000001111111111000000000000000000,
		640'b00000000000000000000000000000000000111111000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001110000111001111111100011110000011110000000000001111000000011100000001110000000000111000011111111100011111110000000000001110000000111111111000000000001111000000001110000111000000000110001100000111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000011111000000000000000000,
		640'b00000000000000000000000000000000000011111110000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001111000010000000001000000000000000100000000000000000000100000000000100000000011111000000111110000000000000000000000001111000000000000000100000000000000000010000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000011110000000000000000000,
		640'b00000000000000000000000000000000000001111111000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000111110000000000000000000,
		640'b00000000000000000000000000000000000000111111100111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000111100000000000000000000,
		640'b00000000000000000000000000000000000000011111111111100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000111100000000000000000000,
		640'b00000000000000000000000000000000000000000111111111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001111111110000000000000000,
		640'b00000000000000000000000000000000000000000011111110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111111110000000000000000,
		640'b00000000000000000000000000000000000000000000111110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000111111110000000000000000,
		640'b00000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000011111110000000000000000,
		640'b00000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000111111100000000000000000,
		640'b00000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111111000000000000000000,
		640'b00000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111111110000000000000000000,
		640'b00000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111111000000000000000000000,
		640'b00000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000,
		640'b00000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000,
		640'b00000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000,
		640'b00000000000000000000000000000011110000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000,
		640'b00000000000000000000000000000111111000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000,
		640'b00000000000000000000000000000111111111000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000,
		640'b00000000000000000000001111000111111111100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000,
		640'b00000000000000000000011111111111111111111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000,
		640'b00000000000000000000011111111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000,
		640'b00000000000000000000001111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000,
		640'b00000000000000000000000111111111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000,
		640'b00000000000000000000000011111111110000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000,
		640'b00000000000000000000000011110000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000,
		640'b00000000000000000000000011110000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000,
		640'b00000000000000000000111111110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000,
		640'b00000000000000000001111111110000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000,
		640'b00000000000000000001111111100000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000,
		640'b00000000000000000001111111100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000,
		640'b00000000000000000001111111110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000,
		640'b00000000000000000000111111111100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000,
		640'b00000000000000000000011111111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000,
		640'b00000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000,
		640'b00000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000,
		640'b00000000000000000000000111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000,
		640'b00000000000011100000000111100011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000,
		640'b00000000000111111110000011100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000,
		640'b00000000000111111111111111110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000,
		640'b00000000000111111111111111110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000,
		640'b00000000000001111111111111100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000,
		640'b00000000000000111111111111100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000,
		640'b00000000000000011111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000,
		640'b00000000000000011111100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000,
		640'b00000000000000001111100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000,
		640'b00000000000000000111100000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000,
		640'b00000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000,
		640'b00000000000000000011110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000,
		640'b00000000000000000111110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000,
		640'b00000000000000001111100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000,
		640'b00000000000000011111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000,
		640'b00000000000011111111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100,
		640'b00000000001111111110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
		640'b00000000001111111000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
		640'b00000000001111110000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110,
		640'b00000000001111111000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000001111100000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,
		640'b00000000000111111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000001111100000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011,
		640'b00000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000111100000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011,
		640'b00000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000111111011111111111111111100000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
		640'b00000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000011111111111100000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011111110000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011111110000000000000000111111111111111111111111100000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000001111100000001111111111111111111111111111111111111111111000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000001111111111110000000000000000000011111111101111111111111000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000001111111111000000000000000000000000000111111000000000000011111111110000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011111111000000000000000000000000000000011111000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000111111110000000000000000000000000000000000111110000000000000000000000000000111111110000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000001111111000000000000000000000000000000000000001111100000000000000000000000000000000011111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111000000000000000000000000000000000000000111110000000000000000000000000000000000000001111110000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110011100001111110000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111110000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000001111110000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000001111110000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000111110000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000001111110000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000111110000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000001111110000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000011111000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000001111100000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000011111000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000011111000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000001111100000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000011111000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000111110000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000011111000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000001111000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000111100000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000011111000000000000000000000000000000000000001111111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001111100000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011110000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001111000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000111100000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001111000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111100000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001110000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111100000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001110000000000000000000000000000000000111110111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111100000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001111000000000000000000000000000000001111110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000011111111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001111000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011110000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001110000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011100000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001110000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111111111111111111111011110000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011100000000000000000000000111111111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000011100000000111111110000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111000000000000000000000011111110000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000011111111000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011110000000000000000000001111110000000011100011110000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000111000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111100000000000000000000111111000000000111000001110000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011100000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111000000000000000000001111110000000001110000001111100000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000011100000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011111000000000000000000111111000000000001110000001111110000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000011110000000000000000000000000000000000001111000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111000000000000000011111100000000000001110000000000111000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000001110000000000000000000000000000000000011111110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001111110000000000000001111110000000000000001100000000000111000000000000000000000000000000000000000000000000000001111000011111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011111110000000000000111111000000000000000001100000000111111000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000011000000000000000000111111100000000001110000001111000000011101111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111101110000000000111111110000000000000000001100000011111111000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000011111111000000000000000000111111000000001111101111111100000011100000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000111001110000000001111110000000000000000000001100000111100000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000011110111100000000000000000000111100000011111111111111110000011100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001110011110000000011110000000000000000000000001100001111000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111000011100000000000000000000111000000011101111110001111000011100000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000011100011100000001111100000000000000000000000001100111100000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000111000011100000000000000000001111000000011000000000000111111011100000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111000011100000111110000000000000000000000000001111111000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000011111001111000011100000000000000000001110000000111000000000000011111111100000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001110000011100001111000000000000000000000000000001111100000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000001111111111110000111000000000000000000011110000000111000000000000000011111000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000011100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111110001111000000000000000000011100000000111000000000000000001111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000011101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000011100000000000011110000000000000000000011100000000111000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000011100000000000111100000000000000000000011100000111110000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000011100000000001111100000000000000000000011111111111100000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000011100000000001111000000000000000000000001111111100000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000011100000000011110000000000000000000000000111110000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000011100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000111100000001111000000001111100000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000001111000000011110000000011111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000111110000000111110000000011011100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000001111111100000000111111111100011111100000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000011111111000000000111111111100011111100000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000111100000000000000000000011100000111000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000111000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000111000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000001111000000000000000000111100000000000000000000000000011111000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000001110000000000000000001110000000000001111110000000000011111100000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000001110000000000000000001110000000000001111111000000000011001110000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000001110000000000000000001110000000000001110111100000000011101110000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000001110000000000000000000000000000000001110000000000000000001110000000000001111011110000000011111111000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000001110000000000000001111110000000000011110000000000000000001110000000000000111100111100000001111110000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000001110000000000000011111111000000000011100000000000000000001110000000000000011110011100000000111100000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000001110000111000000000000000000000000000000000000000000001110111110000000111100111100000000011100000000000000000001110000000000000001111001110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000011100000111000000000000000000000000000000000000000000000111111111100000111000011110000000011100000000111110000001110000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000111000000111100000000000000000000000000000000000000000000111110111111001111000001111111111111100000011111111000001110000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000001111000000111000000011100000000000000000000000000000000000000000000111100000111111110000000111111111111000000111100011100001110000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011111110001110000000011100000000000000000000000000000000000000000000000000000001111000000000001111111100000001111000001110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000011111111001110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000011100111101110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000001111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000011100111111110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000011100011111110000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000001111100011111111000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011111000011110111000000001110000000000000000000000000000000000000000000000000000000000000000011110000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000001111110000111110111000000001110000000000000000000000000000000000000000000000000000000000000000111111000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000001111000000111100111000000001110000000000000000000000000000000000000000000000000000000000000001110111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000001110000001111001110000000000111000000000000000000000000000000000000000000000000000000000000001110011000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000001110000001111001110000000000110000000000000000000000000000000000000000000000000000000000000011110011100000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000001110000001111001110000000000111000000000000000000000000000000000000000000000000000000000000011100011100000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011100000001110001110000000000111000000000000000000111110000000000000000000000000000000000000011100011100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000011100000111110001110000000000111000000000000000001111111000000000000000000000000000000000000011100001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000111100001111100001110000000001110000000000000000011100111000001111100000000000000000000000000011100001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000111111111111000001110000000001110000000000000000111100111000111111110000000000000000000000000111100001110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000001111111111100000001100000000001110000000000000000111000111111111000111000000000000000000000000111000001111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000011111111110000000011100000000000111000000000000001110000011111100000111001110000000000000000000111000000111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000011111100000000000111100000000000111000000000000001110000011110000000111011111110000000000000001111000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011100000000000001111000000000000111000000000000011100000000000000000111111011111111000000000011110000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000011110000000000000011100000000000011100000000000000000111110000011111111110001111100000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000111100000000000000011100000000000111000000000000000000011110000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000001111000000000000000001100000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000001110000000000000000001100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000001110000000000000000011100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000111100000000000000001111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000001111000000000000000011110000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011100000000000000001111000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000011100000000000000011110000000000011100000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000011100000000000001111100000000000011100000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000011000000000000011110000000000000111000000000000000000000000000000000000000000000000000000000000000000001110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000011000000000110111100000000000001111000000000000000000000000000000000000000000000000000000000000000000001110111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000011000000111111111000000000000001110000000000000000000000000000000000000000000000000111111110000000000001110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000011000001111111110000000000000011100000000000000000000000000000000000000000000000111111111111000000000001110001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000011000111110000000000001111111111000000000000000000000000000000000000000000000011111110000111000000000001110000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000011101111100000000000111111111110000000000000000000000000000000000000000000011111100000000011100000000001110000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000011111110000000000001111000000000000000000000000000000000000000000000000000111100000000000011100000000001111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000001111000000000000001100000000000000000000000000000000000000000000000000011110000000000000011100000000000111000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000011110000000000011111100000000000000011100000000000111100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000001111111111111111111110000000000000000011100000000000011110000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000001110111111111111100000000000000000000011100000000000001111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000011110001111100000000000000000000000000011100000000000000111000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000011100000000000000000000000000000000000011100000000000000111100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000111100000000000000000000000000000000000011100000000000000011110000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000001111000000000000000000000000000000000000011110000000000000001111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000011110000000000000000000000000000000000000001110000000000000000111100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000001111100000000000000000000000000000000000000001111000000000000000011100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000111111000000000000000000000111110000000000000000111100000000000000011100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000001111100000000000000000000000111110000000000000000011110000000000000011100000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000011110000000000000000000000001111110000000000000000001111000000000111111100000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000111100000000000000000000000001101111000000000000000000111100000001111111000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000011111000000000000000000000000001100111000000000000000000011110000011111110000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000111100000000000000000000000000001110111000000000000000000001111000011100000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000011111000000000000000000000000000001110111000000000000000000000111100111100000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000111110000000000000000000000000000001110111000000000000000000000011100111100000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000011111000000000000000000000000000000001111111000000000000000000000011100111100000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011111000000000000000000000001111110001111100000000000000000000000000000000000111110000000000000000000000011100011100000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000001111100000000000000000011111111111111111000000000000000000000000000000000000011110000000000000000000000011100011100000000000000000111100000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000011110000000000000011111111111111111100000000000000000000000000000000000000001110000000000000000000000011100011100000000000000000111100000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000111111000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000111100000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011100000000000000000111110000000000000011100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000111111111000000000000000000000000000000000000000111000011100000000000000000011111000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000001111000011100000000000000000001111100000000000111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000001110000001110000000000000000000111110000000000111100000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111111100000000000000011111111111000000000000000000000000011110000001110000000000000000000011111000000000111100000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000011110011111000000000000000000011111111110000000000000000000000000011111110000000000000000000000111100000001110000000000000000000001111000000000111100000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000011100000001111110000000000001111111111100000000000000000000000000000000111111100000000000000000000111000000001110000000000000000000001111000000000111100000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000111100000000011111111111111111111111000000000000000000000000000000000000000111110000000000000000001111000000001110000000000000000000000111000000000111000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000111000000000000111111111111111110000000000000000000000000000000000000000000011111000000000000000001110000000000110000000000000000000000111100000000111000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000001111000000000000000111111001000000000000000000000000000000000000000000000000000111100000000000000011110000000000111000000000000000000000111100000000111100000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000011100111110000111000000000000000000000111100000000111100000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000011111111111100111000000000000000000000011110000000111100000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000011111100011100111000000000000000000000011111000000111000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000100000001110111000000000000000000000001111100000111000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000001111110000000000000000000000000111111111111000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111110000000000000000000000000011111111111000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000000000111111110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000011111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000011111111111101111000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111110000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001111111000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000011111111000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001111000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100001111111111000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111011111100111000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000111000000000000000000000000000000000000000000000000011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000111000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000111100000000000000000000000000000000000000000000000011000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000111111111110000000000000000000000000000000000000000011000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000011000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000001110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000001100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000111000011111111100000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000011100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000001111000000011111110000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000011100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000001111000000000011111100000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000011100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		640'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000001111110000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000011100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

        };

	assign data = ROM[addr];

endmodule