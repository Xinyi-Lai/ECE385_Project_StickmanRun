


//-------------------------------------------------------------------------
//    Star.sv Spring 2020											 --
//    Adapted from Ball.sv, lab8                                         --
//    Real time score keeper on VGA display					             --
//    Indicate how many coins are collected when the player wins.        --
//-------------------------------------------------------------------------

module star ( 	input		Clk,                // 50 MHz clock
							Reset,              // Active-high reset signal
				input [9:0] DrawX, DrawY,       // Current pixel coordinates
				input [2:0] CoinStatus, 	   // Accept from gamelogic
				output logic is_star           // Whether current pixel belongs to star 
 
			  );

	parameter [9:0] Star1_X_Pos = 10'd240; //the rightmost star position
	parameter [9:0] Star1_Y_Pos = 10'd200;  //the leftmost star position

	parameter [9:0] Star2_X_Pos = 10'd300; //the middle star position
	parameter [9:0] Star2_Y_Pos = 10'd200; //the middle star position

	parameter [9:0] Star3_X_Pos = 10'd360;  //the leftmost star position
	parameter [9:0] Star3_Y_Pos = 10'd200;  //the leftmost star position


	parameter [4:0] Star_Height = 5'd16;   // Height of the single score
	parameter [3:0] Star_Width = 4'd8;     // Width of the single score

	logic star_on;         //Tell whether the pixel belongs to star1 or star2 or star3
	
	
	logic [2:0] Collected_Number;           //the number of collected coin

    always_comb begin
		Collected_Number = 3'd0;
		for  (int i=0; i<3; i++) begin
        if ( CoinStatus[i] == 1'b0)
            Collected_Number = Collected_Number + 3'd1;
        else
            Collected_Number = Collected_Number;
		end
    end
	

    //Compute whether the pixel belongs to the score font.
    /* Since the dividers are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are divided. */

	int Scaled_X, Scaled_Y; //the scaled difference betweent th epixel and the origin of score
	
	logic [7:0] sprite_adress;
	logic [0:7] sprite_data;

	always_comb begin

		if ( DrawX >=Star1_X_Pos && DrawX < Star1_X_Pos + Star_Width*5 &&
				DrawY >=Star1_Y_Pos && DrawY < Star1_Y_Pos + Star_Height*5) begin    
			star_on = 1'b1;
			Scaled_X = (DrawX-Star1_X_Pos)/5;
			Scaled_Y = (DrawY-Star1_Y_Pos)/5;
            if (Collected_Number!=3'd0)
			    sprite_adress = Scaled_Y + Star_Height* 8'h1;
            else
                sprite_adress = Scaled_Y + Star_Height* 8'h0;
		end

		else if ( DrawX >=Star2_X_Pos && DrawX < Star2_X_Pos + Star_Width*5 &&
				DrawY >=Star2_Y_Pos && DrawY < Star2_Y_Pos + Star_Height*5) begin    
            star_on = 1'b1;
			Scaled_X = (DrawX-Star2_X_Pos)/5;
			Scaled_Y = (DrawY-Star2_Y_Pos)/5;
            if (Collected_Number==3'd2 || Collected_Number==3'd3)
			    sprite_adress = Scaled_Y + Star_Height* 8'h1;
            else
                sprite_adress = Scaled_Y + Star_Height* 8'h0;
		end
		else if ( DrawX >=Star3_X_Pos && DrawX < Star3_X_Pos + Star_Width*5 &&
				DrawY >=Star3_Y_Pos && DrawY < Star3_Y_Pos + Star_Height*5) begin    
            star_on = 1'b1;
			Scaled_X = (DrawX-Star3_X_Pos)/5;
			Scaled_Y = (DrawY-Star3_Y_Pos)/5;
            if (Collected_Number==3'd3)
			    sprite_adress = Scaled_Y + Star_Height* 8'h1;
            else
                sprite_adress = Scaled_Y + Star_Height* 8'h0;
		end
		else begin
			star_on = 1'b0;
			Scaled_X = 0;
			Scaled_Y = 0;
			sprite_adress = 8'h0;
		end
		

	end

	digits_rom my_digits(.addr(sprite_adress), .data(sprite_data));

	always_comb begin
		if (star_on==1'b1 && sprite_data[Scaled_X]== 1'b1) begin
			is_star = 1'b1;
        end
        else begin
            is_star = 1'b0;
        end
    end

endmodule