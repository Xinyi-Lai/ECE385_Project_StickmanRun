module stickman_rom ( input [10:0] addr, output [83:0] data);

	//parameter ADDR_WIDTH = 11;
	parameter ROM_LENGTH = 120*9;	// 1080
	parameter DATA_WIDTH = 84;
	// logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition: height: 120 * 9, width: 84
	parameter [0:ROM_LENGTH-1][DATA_WIDTH-1:0] ROM = {
		// height: 120, width: 84
		//Page 1
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000001111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000011000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000001111110000000000000000,
		84'b000000000000000000000000000000000000000001111111111111100000001111110000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000011111111000000000000000,
		84'b000000000000000000000000000000000000000011111111111100000000011111111000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000111111111000000000000000,
		84'b000000000000000000000000000000000011111111111111110000000000111111110000000000000000,
		84'b000000000000000000000000000000001111111111111111110000000000111111100000000000000000,
		84'b000000000000000000000000000001111111111111111111111000000001111111100000000000000000,
		84'b000000000000000000000000001111111111111111111111111100000011111111000000000000000000,
		84'b000000000000000000000000111111111111111111111111111100000011111111000000000000000000,
		84'b000000000000000000000001111111111111111111111111111110000011111111000000000000000000,
		84'b000000000000000000000001111111111111111101111111111111000111111110000000000000000000,
		84'b000000000000000000000001111111111111100001111111111111000111111110000000000000000000,
		84'b000000000000000000000001111111111000000001111111111111101111111100000000000000000000,
		84'b000000000000000000000001111111100000000001111111111111111111111100000000000000000000,
		84'b000000000000000000000011111111000000000001111111111111111111111000000000000000000000,
		84'b000000000000000000000011111111000000000001111111111111111111111000000000000000000000,
		84'b000000000000000000000011111111000000000011111111011111111111110000000000000000000000,
		84'b000000000000000000000011111110000000000011111110011111111111110000000000000000000000,
		84'b000000000000000000000011111110000000000011111110001111111111100000000000000000000000,
		84'b000000000000000000000011111110000000000011111110000111111111100000000000000000000000,
		84'b000000000000000000000111111110000000000011111110000111111111100000000000000000000000,
		84'b000000000000000000000111111110000000000011111110000011111111000000000000000000000000,
		84'b000000000000000000000111111110000000000011111110000001111110000000000000000000000000,
		84'b000000000000000000000111111110000000000111111110000001111110000000000000000000000000,
		84'b000000000000000000000111111100000000000111111110000000011100000000000000000000000000,
		84'b000000000000000000000111111100000000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000111111100000000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000111111100000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000001111111100000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000001111111100000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000001111111000000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000001111111000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000001111111000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000001111110000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000111110000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111111111110000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111111111111000000000000000,
		84'b000000000000000000000000000000000000111111110011111111111111111111111100000000000000,
		84'b000000000000000000000000000000000001111111100000011111111111111111111100000000000000,
		84'b000000000000000000000000000000000001111111100000000001111111111111111100000000000000,
		84'b000000000000000000000000000000000011111111000000000000000011111111111100000000000000,
		84'b000000000000000000000000000000000011111111000000000000000000011111111000000000000000,
		84'b000000000000000000000000000000000011111110000000000000000000111111111000000000000000,
		84'b000000000000000000000000000000000111111110000000000000000000111111110000000000000000,
		84'b000000000000000000000000000000000111111110000000000000000001111111110000000000000000,
		84'b000000000000000000000000000000001111111100000000000000000011111111100000000000000000,
		84'b000000000000000000000000000000001111111100000000000000000011111111000000000000000000,
		84'b000000000000000000000000000000001111111000000000000000000111111111000000000000000000,
		84'b000000000000000000000000000000011111111000000000000000000111111110000000000000000000,
		84'b000000000000000000000000000000011111110000000000000000001111111100000000000000000000,
		84'b000000000000000000000000000000111111110000000000000000011111111100000000000000000000,
		84'b000000000000000000000000000000111111110000000000000000011111111000000000000000000000,
		84'b000000000000000000000000000001111111100000000000000000111111111000000000000000000000,
		84'b000000000000000000000000000001111111100000000000000001111111110000000000000000000000,
		84'b000000000000000000000000000011111111000000000000000001111111100000000000000000000000,
		84'b000000000000000000000000000111111111000000000000000011111111100000000000000000000000,
		84'b000000000000000000000000001111111111000000000000000011111111000000000000000000000000,
		84'b000000000000000000000000011111111110000000000000000111111111000000000000000000000000,
		84'b000000000000000000000001111111111110000000000000001111111110000000000000000000000000,
		84'b000000000000000000000011111111111100000000000000001111111100000000000000000000000000,
		84'b000000000000000000000111111111111000000000000000011111111100000000000000000000000000,
		84'b000000000000000000001111111111110000000000000000011111111110000000000000000000000000,
		84'b000000000000000000111111111111000000000000000000001111111111000000000000000000000000,
		84'b000000000000000000111111111110000000000000000000001111111111000000000000000000000000,
		84'b000000000000000011111111111100000000000000000000000111111111100000000000000000000000,
		84'b000000000000000111111111110000000000000000000000000001111111000000000000000000000000,
		84'b000000000000001111111111100000000000000000000000000000111111000000000000000000000000,
		84'b000000000000011111111111000000000000000000000000000000011110000000000000000000000000,
		84'b000000000001111111111110000000000000000000000000000000000000000000000000000000000000,
		84'b000000000011111111111000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000111111111110000000000000000000000000000000000000000000000000000000000000000,
		84'b000000001111111111100000000000000000000000000000000000000000000000000000000000000000,
		84'b000000001111111111000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000001111111110000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000001111111100000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000001111111100000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000111111100000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000111111100000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000111111110000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000011111100000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000011111000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

		//Page 2
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000011111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000110000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100011111000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100011111100000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100111111100000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000111111100000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000111111100000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000111111100000000000000000,
		84'b000000000000000000000000000000000000000000111111111111100000111111100000000000000000,
		84'b000000000000000000000000000000000000000000111111111110000001111111100000000000000000,
		84'b000000000000000000000000000000000000000111111111110000000001111111000000000000000000,
		84'b000000000000000000000000000000000000011111111111110000000001111111000000000000000000,
		84'b000000000000000000000000000000000011111111111111111000000001111111000000000000000000,
		84'b000000000000000000000000000000000111111111111111111100000011111111000000000000000000,
		84'b000000000000000000000000000000111111111111111111111110000011111111000000000000000000,
		84'b000000000000000000000000000111111111111111111111111111100011111111000000000000000000,
		84'b000000000000000000000000011111111111111111111111111111100011111110000000000000000000,
		84'b000000000000000000000000111111111111111111111111111111110011111110000000000000000000,
		84'b000000000000000000000000111111111111111001111111111111111111111110000000000000000000,
		84'b000000000000000000000000111111111111100001111111111111111111111110000000000000000000,
		84'b000000000000000000000001111111111100000001111111011111111111111100000000000000000000,
		84'b000000000000000000000001111111110000000001111111001111111111111100000000000000000000,
		84'b000000000000000000000001111111000000000001111111000111111111111100000000000000000000,
		84'b000000000000000000000001111111000000000011111111000011111111111100000000000000000000,
		84'b000000000000000000000001111111000000000011111111000001111111111100000000000000000000,
		84'b000000000000000000000001111111000000000011111111000000111111111000000000000000000000,
		84'b000000000000000000000001111111000000000011111110000000001111111000000000000000000000,
		84'b000000000000000000000001111111000000000011111110000000001111111000000000000000000000,
		84'b000000000000000000000011111111000000000011111110000000000111110000000000000000000000,
		84'b000000000000000000000011111111000000000011111110000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000000011111110000000000000000000000000000000000000,
		84'b000000000000000000000011111110000000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111110000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111110000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000111111110000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000111111110000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000111111110000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000111111110000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000111111110000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000111111100000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111100000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000001111000000000001111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111111110000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111111111111111111000000000000000,
		84'b000000000000000000000000000000000011111111101111111111111111111111111100000000000000,
		84'b000000000000000000000000000000000011111111000001111111111111111111111100000000000000,
		84'b000000000000000000000000000000000111111111000000000011111111111111111100000000000000,
		84'b000000000000000000000000000000001111111110000000000000011111111111111100000000000000,
		84'b000000000000000000000000000000001111111100000000000000000000111111111100000000000000,
		84'b000000000000000000000000000000011111111100000000000000000000000111111100000000000000,
		84'b000000000000000000000000000000111111111000000000000000000000001111111100000000000000,
		84'b000000000000000000000000000000111111110000000000000000000000001111111100000000000000,
		84'b000000000000000000000000000001111111110000000000000000000000001111111000000000000000,
		84'b000000000000000000000000000011111111100000000000000000000000001111111000000000000000,
		84'b000000000000000000000000000011111111100000000000000000000000001111111000000000000000,
		84'b000000000000000000000000000111111111000000000000000000000000011111111000000000000000,
		84'b000000000000000000000000001111111110000000000000000000000000011111111000000000000000,
		84'b000000000000000000000000001111111100000000000000000000000000011111111000000000000000,
		84'b000000000000000000000000011111111100000000000000000000000000011111110000000000000000,
		84'b000000000000000000000000111111111000000000000000000000000000011111110000000000000000,
		84'b000000000000000000000001111111111000000000000000000000000000011111110000000000000000,
		84'b000000000000000000000111111111110000000000000000000000000000011111110000000000000000,
		84'b000000000000000000001111111111100000000000000000000000000000111111110000000000000000,
		84'b000000000000000000111111111111000000000000000000000000000000111111110000000000000000,
		84'b000000000000000001111111111111000000000000000000000000000000111111100000000000000000,
		84'b000000000000000011111111111100000000000000000000000000000000111111100000000000000000,
		84'b000000000000001111111111111000000000000000000000000000000000111111100000000000000000,
		84'b000000000000011111111111100000000000000000000000000000000001111111100000000000000000,
		84'b000000000000111111111111000000000000000000000000000000000001111111100000000000000000,
		84'b000000000011111111111110000000000000000000000000000000000001111111100000000000000000,
		84'b000000001111111111111000000000000000000000000000000000000001111111100000000000000000,
		84'b000000011111111111110000000000000000000000000000000000000001111111111000000000000000,
		84'b000000111111111111000000000000000000000000000000000000000001111111111000000000000000,
		84'b000011111111111110000000000000000000000000000000000000000001111111111100000000000000,
		84'b000111111111111000000000000000000000000000000000000000000000111111111100000000000000,
		84'b000111111111110000000000000000000000000000000000000000000000011111111100000000000000,
		84'b001111111111100000000000000000000000000000000000000000000000000111111100000000000000,
		84'b001111111110000000000000000000000000000000000000000000000000000011111000000000000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000011111100000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000011111100000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000001111000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

		//Page 3
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000001111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111111000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110111111100000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111100111111100000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000111111100000000000000000000,
		84'b000000000000000000000000000000000000000001111111111100000111111100000000000000000000,
		84'b000000000000000000000000000000000000000111111111110000000111111100000000000000000000,
		84'b000000000000000000000000000000000000001111111111111000000111111100000000000000000000,
		84'b000000000000000000000000000000000000111111111111111100000111111100000000000000000000,
		84'b000000000000000000000000000000000011111111111111111110000111111100000000000000000000,
		84'b000000000000000000000000000000001111111111111111111111100111111100000000000000000000,
		84'b000000000000000000000000000000111111111111111111111111110111111100000000000000000000,
		84'b000000000000000000000000000011111111111111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000111111111111111111111111111111111111100000000000000000000,
		84'b000000000000000000000000011111111111111101111111111111111111111100000000000000000000,
		84'b000000000000000000000000011111111111110001111111011111111111111100000000000000000000,
		84'b000000000000000000000000111111111111000001111111001111111111111100000000000000000000,
		84'b000000000000000000000000111111111100000001111111000011111111111100000000000000000000,
		84'b000000000000000000000000111111111000000001111111000001111111111100000000000000000000,
		84'b000000000000000000000000011111110000000011111111000000111111111100000000000000000000,
		84'b000000000000000000000000011111110000000011111111000000011111111100000000000000000000,
		84'b000000000000000000000000011111110000000011111110000000000111111100000000000000000000,
		84'b000000000000000000000000011111110000000011111110000000000011111000000000000000000000,
		84'b000000000000000000000000011111110000000011111110000000000001110000000000000000000000,
		84'b000000000000000000000000011111110000000011111110000000000000000000000000000000000000,
		84'b000000000000000000000000011111110000000011111110000000000000000000000000000000000000,
		84'b000000000000000000000000011111110000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000000011111110000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000000011111110000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000000111111110000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111000001111111110000000000000000000000000000000000000,
		84'b000000000000000000000000001111110000001111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000111100000001111111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000000000000111111110111111111111111111111111000000000000000,
		84'b000000000000000000000000000000000000111111100001111111111111111111111000000000000000,
		84'b000000000000000000000000000000000001111111100000000111111111111111111100000000000000,
		84'b000000000000000000000000000000000001111111100000000000111111111111111100000000000000,
		84'b000000000000000000000000000000000001111111000000000000000011111111111100000000000000,
		84'b000000000000000000000000000000000011111111000000000000000000011111111100000000000000,
		84'b000000000000000000000000000000000011111111000000000000000000000111111100000000000000,
		84'b000000000000000000000000000000000011111110000000000000000000000111111100000000000000,
		84'b000000000000000000000000000000000111111110000000000000000000000111111110000000000000,
		84'b000000000000000000000000000000000111111110000000000000000000000111111110000000000000,
		84'b000000000000000000000000000000000111111100000000000000000000000011111110000000000000,
		84'b000000000000000000000000000000001111111100000000000000000000000011111110000000000000,
		84'b000000000000000000000000000000001111111100000000000000000000000011111110000000000000,
		84'b000000000000000000000000000000001111111000000000000000000000000011111110000000000000,
		84'b000000000000000000000000000000011111111000000000000000000000000011111111000000000000,
		84'b000000000000000000000000000000011111111000000000000000000000000011111111000000000000,
		84'b000000000000000000000000000000111111110000000000000000000000000001111111000000000000,
		84'b000000000000000000000000000101111111110000000000000000000000000001111111000000000000,
		84'b000000000000000000000111111111111111110000000000000000000000000001111111000000000000,
		84'b000000000000000111111111111111111111100000000000000000000000000001111111000000000000,
		84'b000000000111111111111111111111111111100000000000000000000000000001111111100000000000,
		84'b000001111111111111111111111111111111100000000000000000000000000001111111100000000000,
		84'b000011111111111111111111111111111111000000000000000000000000000001111111100000000000,
		84'b000011111111111111111111111111111110000000000000000000000000000001111111100000000000,
		84'b000011111111111111111111111111100000000000000000000000000000000000111111100000000000,
		84'b000111111111111111111111100000000000000000000000000000000000000000111111100000000000,
		84'b000111111111111111000000000000000000000000000000000000000000000000111111111100000000,
		84'b000111111111000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000111111100000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000111111000000000000000000000000000000000000000000000000000000000011111111111000000,
		84'b000001100000000000000000000000000000000000000000000000000000000000000111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

		//Page 4
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000001111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111111111000000000000001111110000000000000,
		84'b000000000000000000000000000000111111111111111111111000000000001111111111000000000000,
		84'b000000000000000000000000000001111111111011111111111100000011111111111111000000000000,
		84'b000000000000000000000000000001111111110011111111111100011111111111111111000000000000,
		84'b000000000000000000000000000001111111100011111111111111111111111111111111000000000000,
		84'b000000000000000000000000000001111111000011111111111111111111111111111111000000000000,
		84'b000000000000000000000000000001111111000011111111111111111111111111111110000000000000,
		84'b000000000000000000000000000001111111000011111111111111111111111111110000000000000000,
		84'b000000000000000000000000000001111111100111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000111111100111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000111111100111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000111111100111111101111111000000000000000000000000000000,
		84'b000000000000000000000000000000111111100111111100010000000000000000000000000000000000,
		84'b000000000000000000000000000000111111100111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111110111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111110111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000011111110111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000111111110011111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000111111110001111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000111111110000111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000111111100000011111111111000000000000000000000000,
		84'b000000000000000000000000000000000000111111100000001111111111100000000000000000000000,
		84'b000000000000000000000000000000000000111111100000000011111111110000000000000000000000,
		84'b000000000000000000000000000000000001111111100000000001111111111000000000000000000000,
		84'b000000000000000000000000000000000001111111100000000000111111111100000000000000000000,
		84'b000000000000000000000000000000000001111111100000000000011111111110000000000000000000,
		84'b000000000011111000000000000000000001111111000000000000001111111110000000000000000000,
		84'b000000000111111111110000000000000001111111000000000000000111111110000000000000000000,
		84'b000000001111111111111111100000000001111111000000000000000011111111000000000000000000,
		84'b000000011111111111111111111111100001111111000000000000000011111111000000000000000000,
		84'b000000111111111111111111111111111111111111000000000000000001111111000000000000000000,
		84'b000001111111111111111111111111111111111111000000000000000001111111100000000000000000,
		84'b000001111111111111111111111111111111111111000000000000000001111111100000000000000000,
		84'b000001111111111111111111111111111111111110000000000000000000111111110000000000000000,
		84'b000001111111000000111111111111111111111110000000000000000000111111110000000000000000,
		84'b000000111110000000000011111111111111111110000000000000000000011111110000000000000000,
		84'b000000011100000000000000000011111111111110000000000000000000011111111000000000000000,
		84'b000000000000000000000000000000000111111100000000000000000000011111111000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000001111111000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000001111111100000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111100000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111110000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111110000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000011111110000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000011111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000011111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000001111111100000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000001111111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000111111111111000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000011111111111000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000011111111111000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000001111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

		//Page 5
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000011111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000001111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111111000000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111111100000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111111100000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000000000000011111111100000011111111111111000000000000000000,
		84'b000000000000000000000000000000000000011111111100000000000000111110000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111101111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100011111111111000000000000000000000000,
		84'b000000000000011111111000000000000000000111111100001111111111100000000000000000000000,
		84'b000000000000111111111110000000000000000111111100000111111111100000000000000000000000,
		84'b000000000001111111111111110000000000000111111100000011111111110000000000000000000000,
		84'b000000000011111111111111111110000000000111111100000001111111111000000000000000000000,
		84'b000000000011111111111111111111100000000111111100000000111111111100000000000000000000,
		84'b000000000001111111111111111111111000000111111100000000011111111100000000000000000000,
		84'b000000000001111111111111111111111111000111111100000000001111111100000000000000000000,
		84'b000000000000011111011111111111111111110111111100000000000111111110000000000000000000,
		84'b000000000000000000000111111111111111111111111100000000000111111110000000000000000000,
		84'b000000000000000000000000111111111111111111111100000000000011111111000000000000000000,
		84'b000000000000000000000000001111111111111111111100000000000011111111000000000000000000,
		84'b000000000000000000000000000001111111111111111100000000000011111111000000000000000000,
		84'b000000000000000000000000000000011111111111111100000000000001111111100000000000000000,
		84'b000000000000000000000000000000000011111111111110000000000001111111100000000000000000,
		84'b000000000000000000000000000000000000111111111100000000000000111111100000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000111111110000000000000000,
		84'b000000000000000000000000000000000000000001110000000000000000111111110000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000011111111000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000011111111000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000001111111000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000001111111100000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000001111111100000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111100000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111110000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111110000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000011111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000011111111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000001111111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000001111111111111000000,
		84'b000000000000000000000000000000000000000000000000000000000000000001111111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000111111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000111111111110000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000011111111000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

		//Page 6
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000011111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000001111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000001111111101111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111100100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111000000000000000000000000000000,
		84'b000000000000000000111111110000000000000001111111111111100000000000000000000000000000,
		84'b000000000000000001111111111100000000000001111111111111100000000000000000000000000000,
		84'b000000000000000011111111111111100000000001111111111111110000000000000000000000000000,
		84'b000000000000000011111111111111111000000001111111111111111000000000000000000000000000,
		84'b000000000000000011111111111111111110000001111111111111111000000000000000000000000000,
		84'b000000000000000011111111111111111111100000111111111111111100000000000000000000000000,
		84'b000000000000000001111111111111111111111000111111101111111110000000000000000000000000,
		84'b000000000000000000101000111111111111111110111111111111111111000000000000000000000000,
		84'b000000000000000000000000001111111111111111111111110111111111000000000000000000000000,
		84'b000000000000000000000000000011111111111111111111110011111111000000000000000000000000,
		84'b000000000000000000000000000000111111111111111111110001111111100000000000000000000000,
		84'b000000000000000000000000000000000111111111111111111001111111100000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111000111111100000000000000000000000,
		84'b000000000000000000000000000000000000111111111111111000111111110000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111000111111110000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111000011111110000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111000011111111000000000000000000000,
		84'b000000000000000000000000000000000000000000000111110000011111111000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000001111111000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000001111111000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000001111111100000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000001111111100000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000111111100000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000111111110000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000011111110000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000011111111000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000011111111000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000011111111000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000001111111000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000001111111100000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000001111111100000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000001111111111100000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000111111111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000111111111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000111111111111100000000000,
		84'b000000000000000000000000000000000000000000000000000000000000011111111111100000000000,
		84'b000000000000000000000000000000000000000000000000000000000000011111111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000001111111111000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000111111000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,

		//Page 7
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111111111111000000000000000000000,
		84'b000000000000000000000000000000000001111111111101111111111111111111000000000000000000,
		84'b000000000000000000000000000000000001111111111100011111111111111111100000000000000000,
		84'b000000000000000000000000000000000001111111111100000111111111111111110000000000000000,
		84'b000000000000000000000000000000000001111111111100000000111111111111110000000000000000,
		84'b000000000000000000000000000000000000111111111100000000001111111111110000000000000000,
		84'b000000000000000000000000000000000000111111111100000000000001111111100000000000000000,
		84'b000000000000000000000000000000000000111111111000000000000000011111000000000000000000,
		84'b000000000000000000000000000000000000111111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111110000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111110000000000000000000000000000000,
		84'b000000000000000000000000000011000000000001111111111111000000000000000000000000000000,
		84'b000000000000000000000000000111111111000001111111111111000000000000000000000000000000,
		84'b000000000000000000000000001111111111111001111111111111100000000000000000000000000000,
		84'b000000000000000000000000111111111111111111111111111111110000000000000000000000000000,
		84'b000000000000000000000001111111111111111111111111111111110000000000000000000000000000,
		84'b000000000000000000000011111111111111111111111111111111111000000000000000000000000000,
		84'b000000000000000000000011111111111111111111111111111111111100000000000000000000000000,
		84'b000000000000000000000011111111111111111111111111111111111100000000000000000000000000,
		84'b000000000000000000000011111111000111111111111111111111111100000000000000000000000000,
		84'b000000000000000000000001111110000000011111111111111111111100000000000000000000000000,
		84'b000000000000000000000000011000000000000000111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111011111000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111000000000000000000000000000000000,

		//Page 8
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000011111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111110000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111110000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111111111111100000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111111111111100000000000000011111000000000000000,
		84'b000000000000000000000000000000111111111111111111110000000000111111111000000000000000,
		84'b000000000000000000000000000001111111111011111111110000001111111111111100000000000000,
		84'b000000000000000000000000000001111111110011111111110011111111111111111100000000000000,
		84'b000000000000000000000000000001111111100011111111111111111111111111111100000000000000,
		84'b000000000000000000000000000011111111000011111111111111111111111111111000000000000000,
		84'b000000000000000000000000000011111111000011111111111111111111111111111000000000000000,
		84'b000000000000000000000000000011111111000111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000011111110000111111111111111111111111000000000000000000000,
		84'b000000000000000000000000000111111110000111111111111111111110000000000000000000000000,
		84'b000000000000000000000000000111111110000111111111111111100000000000000000000000000000,
		84'b000000000000000000000000000111111100000111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000111111100000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111100000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111100000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111100000111111100000000000000000000000000000000000000,
		84'b000000000000000000000000001111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000011111111000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000011111110000001111111000000000000000000000000000000000000000,
		84'b000000000000000000000000011111110000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000111111110000001111111110000000000000000000000000000000000000,
		84'b000000000000000000000000111111110000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000000111111100000001111111111110000000000000000000000000000000000,
		84'b000000000000000000000000111111100000001111111111111100000000000000000000000000000000,
		84'b000000000000000000000000111111100000001111111111111110000000000000000000000000000000,
		84'b000000000000000000000000011111000000001111111111111111100000000000000000000000000000,
		84'b000000000000000000000000001110000000001111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000001111111100011111111111110000000000000000000000,
		84'b000000000000000000000000000000000000001111111100001111111111111100000000000000000000,
		84'b000000000000000000000000000000000000001111111100000011111111111111000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000111111111111000000000000000000,
		84'b000000000000000000000000000000000000001111111100111111111111111111100000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111111111100000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111111111100000000000000000,
		84'b000000000000000000000000000000000001111111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111111111111110000000000000000000,
		84'b000000000000000000000000000000000011111111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000011111111111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111111000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000011111110000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111110000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000111111110000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111100000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111100000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000111111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111100000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111100000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000011111111100000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111111000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111111000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000001111111110000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000,

		//Page 9
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000001111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000000111111111111111111000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000000000111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000000000001111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000000000011111111100000000000000000000110000000000000,
		84'b000000000000000000000000000000000000001111111111100000000000000000011111000000000000,
		84'b000000000000000000000000000000000000111111111111110000000000000000111111100000000000,
		84'b000000000000000000000000000000000001111111111111110000000000000001111111100000000000,
		84'b000000000000000000000000000000000111111111111111111000000000000011111111100000000000,
		84'b000000000000000000000000000000011111111111111111111100000000000111111111100000000000,
		84'b000000000000000000000000000001111111111111111111111100000000001111111111000000000000,
		84'b000000000000000000000000000111111111111111111111111110000000011111111110000000000000,
		84'b000000000000000000000000001111111111111111111111111110000000111111111100000000000000,
		84'b000000000000000000000000011111111111111001111111111111000001111111111000000000000000,
		84'b000000000000000000000000011111111111100001111111111111000011111111110000000000000000,
		84'b000000000000000000000000011111111110000001111111111111100111111111100000000000000000,
		84'b000000000000000000000000111111111000000011111111111111101111111111000000000000000000,
		84'b000000000000000000000000111111100000000011111111111111111111111110000000000000000000,
		84'b000000000000000000000000111111100000000011111110111111111111111100000000000000000000,
		84'b000000000000000000000000111111100000000011111110011111111111111000000000000000000000,
		84'b000000000000000000000000111111100000000011111110011111111111110000000000000000000000,
		84'b000000000000000000000000111111100000000011111110001111111111110000000000000000000000,
		84'b000000000000000000000000111111100000000011111110000111111111000000000000000000000000,
		84'b000000000000000000000000111111100000000011111110000111111110000000000000000000000000,
		84'b000000000000000000000001111111100000000111111110000011111110000000000000000000000000,
		84'b000000000000000000000001111111100000000111111110000011111100000000000000000000000000,
		84'b000000000000000000000001111111000000000111111110000000110000000000000000000000000000,
		84'b000000000000000000000001111111000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000001111111000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000001111111000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000001111111000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000001111111000000000111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000011111110000000001111111100000000000000000000000000000000000000,
		84'b000000000000000000000001111110000000001111111111100000000000000000000000000000000000,
		84'b000000000000000000000001111100000000001111111111111100000000000000000000000000000000,
		84'b000000000000000000000000011000000000001111111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000001111111111111111111111100000000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111100000000000000000000,
		84'b000000000000000000000000000000000000011111111111111111111111111111000000000000000000,
		84'b000000000000000000000000000000000000011111111011111111111111111111110000000000000000,
		84'b000000000000000000000000000000000000011111110000001111111111111111111000000000000000,
		84'b000000000000000000000000000000000000011111110000000001111111111111111000000000000000,
		84'b000000000000000000000000000000000000011111110000000000001111111111111000000000000000,
		84'b000000000000000000000000000000000000011111110000000000000011111111111000000000000000,
		84'b000000000000000000000000000000000000011111110000000000000111111111111000000000000000,
		84'b000000000000000000000000000000000000011111110000000000001111111111110000000000000000,
		84'b000000000000000000000000000000000000011111110000000000111111111111000000000000000000,
		84'b000000000000000000000000000000000000111111110000000001111111111110000000000000000000,
		84'b000000000000000000000000000000000000111111110000000011111111111100000000000000000000,
		84'b000000000000000000000000000000000000111111110000000111111111111000000000000000000000,
		84'b000000000000000000000000000000000000111111100000011111111111100000000000000000000000,
		84'b000000000000000000000000000000000000111111100000111111111111000000000000000000000000,
		84'b000000000000000000000000000000000000111111100001111111111110000000000000000000000000,
		84'b000000000000000000000000000000000000111111100111111111111100000000000000000000000000,
		84'b000000000000000000000000000000000000111111101111111111110000000000000000000000000000,
		84'b000000000000000000000000000000000000111111111111111111100000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111111000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000001111111111111111000000000000000000000000000000000,
		84'b000000000000000000000000000000000011111111111111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111011111111100000000000000000000000000000000,
		84'b000000000000000000000000000000000111111111001111111100000000000000000000000000000000,
		84'b000000000000000000000000000000001111111110001111111100000000000000000000000000000000,
		84'b000000000000000000000000000000011111111110000111111100000000000000000000000000000000,
		84'b000000000000000000000000000000111111111100000011111000000000000000000000000000000000,
		84'b000000000000000000000000000000111111111000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000001111111110000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000011111111100000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000111111111000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000001111111110000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000001111111110000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000011111111100000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000111111111000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000001111111110000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000011111111110000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000111111111100000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000111111111000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000001111111111000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000011111111100000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000011111111100000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000011111111100000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000011111111110000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000011111111111000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000111111111000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000011111111000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000001111110000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000111100000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000

        };

	assign data = ROM[addr];

endmodule  