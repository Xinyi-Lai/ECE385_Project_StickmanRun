//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf 03-01-2006                               --
//                              03-12-2007                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  12-08-2017                               --
//    Spring 2018 Distribution                                           --
//                                                                       --
//    For use with ECE 385 Lab 8                                         --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------


module  ball (  input         Clk,                // 50 MHz clock
                             Reset,              // Active-high reset signal
                             frame_clk,          // The clock indicating a new frame (~60Hz)
				input [7:0]   keycode, 				 // Accept the last received key 
                input [9:0]   DrawX, DrawY,       // Current pixel coordinates
                output logic  is_ball,             // Whether current pixel belongs to ball or background
			    output logic  is_black
				
				  );
    
    parameter [9:0] Ball_X_Center = 10'd28;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center = 10'd28;  // Center position on the Y axis
    // parameter [9:0] Ball_X_Min = 10'd0;       // Leftmost point on the X axis
    // parameter [9:0] Ball_X_Max = 10'd639;     // Rightmost point on the X axis
    // parameter [9:0] Ball_Y_Min = 10'd0;       // Topmost point on the Y axis
    // parameter [9:0] Ball_Y_Max = 10'd479;     // Bottommost point on the Y axis
    // parameter [9:0] Ball_X_Step = 10'd1;      // Step size on the X axis
    // parameter [9:0] Ball_Y_Step = 10'd1;      // Step size on the Y axis
    parameter [9:0] Ball_Size = 10'd8;        // Ball size
    parameter [16:0] frame_counter_max =16'd2047 ;
	 
	parameter [9:0] earth_height = 10'd20; 	 //Define the earth line
    parameter [9:0] obstacle_height = 10'd40; 
    parameter [9:0] pitfall_height = 10'd00; 
	parameter [9:0] Screen_max = 10'd639;     // Rightmost point on the X axis of the screen

    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
    logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
    logic [15:0] frame_counter;
    logic [9:0] height[frame_counter_max+Screen_max];

    

    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    // Update registers
    always_ff @ (posedge Clk)
    begin
        if (Reset)
        begin
            Ball_X_Pos <= Ball_X_Center;
            Ball_Y_Pos <= Ball_Y_Center;
            Ball_X_Motion <= 10'd0;
            Ball_Y_Motion <= 10'd0;
            frame_counter <= 16'd0;
        end
        else
        begin
            Ball_X_Pos <= Ball_X_Pos_in;
            Ball_Y_Pos <= Ball_Y_Pos_in;
            Ball_X_Motion <= Ball_X_Motion_in;
            Ball_Y_Motion <= Ball_Y_Motion_in;
            
        end
    end
    //////// Do not modify the always_ff blocks. ////////
    always_comb
    begin
        for (int i=0; i<300; i++) begin
			height[i] = earth_height;
		end

        for (int i=300; i<40; i++) begin
            height[i] = pitfall_height;
        end

        for (int i=340; i<800;i++) begin
            height[i] = earth_height;
        end

        for (int i=800; i<840;i++) begin
            height[i] = obstacle_height;
        end

        for (int i=840; i<frame_counter_max+Screen_max;i++) begin
            height[i] = earth_height;
        end
        
    end
    // You need to modify always_comb block.
    always_comb
    begin
        // By default, keep motion and position unchanged
        Ball_X_Pos_in = Ball_X_Pos;
        Ball_Y_Pos_in = Ball_Y_Pos;
        Ball_X_Motion_in = Ball_X_Motion;
        Ball_Y_Motion_in = Ball_Y_Motion;
        
        // Update position and motion only at rising edge of frame clock
        if (frame_clk_rising_edge)
        begin

            Ball_X_Motion_in = 10'd0;
            Ball_Y_Motion_in = 10'd0;
            if (frame_counter<=frame_counter_max)
                frame_counter <= frame_counter+1;
            else 
                frame_counter <= frame_counter_max;
            // Be careful when using comparators with "logic" datatype because compiler treats 
            //   both sides of the operator as UNSIGNED numbers.
            // e.g. Ball_Y_Pos - Ball_Size <= Ball_Y_Min 
            // If Ball_Y_Pos is 0, then Ball_Y_Pos - Ball_Size will not be -4, but rather a large positive number.
            // if( Ball_Y_Pos + Ball_Size >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
			// 		begin
			// 			Ball_X_Motion_in = 10'd0; 
			// 			Ball_Y_Motion_in = (~(Ball_Y_Step) + 1'b1);  // 2's complement.
			// 		end
            // else if ( Ball_Y_Pos <= Ball_Y_Min + Ball_Size )  // Ball is at the top edge, BOUNCE!
			// 		begin
			// 		 Ball_Y_Motion_in = Ball_Y_Step;
			// 		 Ball_X_Motion_in = 10'd0;
			// 		end
            // // TODO: Add other boundary detections and handle keypress here.
			// 	// X boundary detection
            // else if( Ball_X_Pos + Ball_Size >= Ball_X_Max )  // Ball is at the right edge, BOUNCE!
            //    begin
			// 		 Ball_X_Motion_in = (~(Ball_X_Step) + 1'b1);  // 2's complement.
			// 		 Ball_Y_Motion_in = 10'd0; 
			// 		end
            // else if ( Ball_X_Pos <= Ball_X_Min + Ball_Size )  // Ball is at the left edge, BOUNCE!
            //    begin
			// 		 Ball_X_Motion_in = Ball_X_Step; 
			// 		 Ball_Y_Motion_in = 10'd0; 
			// 		end 
			// 	//handle keypress
			// 	else
			// 		begin
			// 			unique case (keycode)
			// 				//press "A", direction is left
			// 				8'h04:
			// 				begin
			// 					Ball_X_Motion_in = (~(Ball_X_Step) + 1'b1); 
			// 					Ball_Y_Motion_in = 10'd0; 
			// 				end	
			// 				//press "D", direction is right
			// 				8'h07:
			// 				begin
			// 					Ball_X_Motion_in = Ball_X_Step; 
			// 					Ball_Y_Motion_in = 10'd0; 
			// 				end
			// 				//press "S", direction is down
			// 				8'h16:
			// 				begin
			// 					Ball_X_Motion_in = 10'd0; 
			// 					Ball_Y_Motion_in = Ball_Y_Step; 
			// 				end
			// 				//press "W", direction is up
			// 				8'h1a:
			// 				begin
			// 					Ball_X_Motion_in = 10'd0; 
			// 					Ball_Y_Motion_in = (~(Ball_Y_Step) + 1'b1); 
			// 				end

			// 				// the key is not pressed, or is released, the key code will be 0x00 (No Event)
			// 				8'h00:
			// 				begin
			// 					Ball_X_Motion_in = Ball_X_Motion; 
			// 					Ball_Y_Motion_in = Ball_Y_Motion; 
			// 				end
			// 				default: ;
			// 			endcase
			// 		end
            // Update the ball's position with its motion
            Ball_X_Pos_in = Ball_X_Pos + Ball_X_Motion;
            Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;
        end
        
        /**************************************************************************************
            ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
            Hidden Question #2/2:
               Notice that Ball_Y_Pos is updated using Ball_Y_Motion. 
              Will the new value of Ball_Y_Motion be used when Ball_Y_Pos is updated, or the old? 
              What is the difference between writing
                "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;" and 
                "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion_in;"?
              How will this impact behavior of the ball during a bounce, and how might that interact with a response to a keypress?
              Give an answer in your Post-Lab.
        **************************************************************************************/
    end
    
    // Compute whether the pixel corresponds to ball or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
    int DistX, DistY, Size;
    assign DistX = DrawX - Ball_X_Pos;
    assign DistY = DrawY - Ball_Y_Pos;
    assign Size = Ball_Size;
    always_comb begin

    //Judge whether the pixel is black
        if (DrawY<=height[frame_counter+DrawX]) //get the height threshold  
            is_black = 1'b1;
        else
            is_black = 1'b0;

        if ( ( DistX*DistX + DistY*DistY) <= (Size*Size) ) 
            is_ball = 1'b1;
        else
            is_ball = 1'b0;
        /* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while 
           the single line is quite powerful descriptively, it causes the synthesis tool to use up three
           of the 12 available multipliers on the chip! */
    end
    
endmodule
